
module openMSP430(aclk, aclk_en, dbg_freeze, dbg_i2c_sda_out, dbg_uart_txd, dco_enable, dco_wkup, dmem_addr_0_, dmem_addr_1_, dmem_addr_2_, dmem_addr_3_, dmem_addr_4_, dmem_addr_5_, dmem_addr_6_, dmem_addr_7_, dmem_addr_8_, dmem_addr_9_, dmem_addr_10_, dmem_addr_11_, dmem_addr_12_, dmem_cen, dmem_din_0_, dmem_din_1_, dmem_din_2_, dmem_din_3_, dmem_din_4_, dmem_din_5_, dmem_din_6_, dmem_din_7_, dmem_din_8_, dmem_din_9_, dmem_din_10_, dmem_din_11_, dmem_din_12_, dmem_din_13_, dmem_din_14_, dmem_din_15_, dmem_wen_0_, dmem_wen_1_, irq_acc_0_, irq_acc_1_, irq_acc_2_, irq_acc_3_, irq_acc_4_, irq_acc_5_, irq_acc_6_, irq_acc_7_, irq_acc_8_, irq_acc_9_, irq_acc_10_, irq_acc_11_, irq_acc_12_, irq_acc_13_, lfxt_enable, lfxt_wkup, mclk, dma_dout_0_, dma_dout_1_, dma_dout_2_, dma_dout_3_, dma_dout_4_, dma_dout_5_, dma_dout_6_, dma_dout_7_, dma_dout_8_, dma_dout_9_, dma_dout_10_, dma_dout_11_, dma_dout_12_, dma_dout_13_, dma_dout_14_, dma_dout_15_, dma_ready, dma_resp, per_addr_0_, per_addr_1_, per_addr_2_, per_addr_3_, per_addr_4_, per_addr_5_, per_addr_6_, per_addr_7_, per_addr_8_, per_addr_9_, per_addr_10_, per_addr_11_, per_addr_12_, per_addr_13_, per_din_0_, per_din_1_, per_din_2_, per_din_3_, per_din_4_, per_din_5_, per_din_6_, per_din_7_, per_din_8_, per_din_9_, per_din_10_, per_din_11_, per_din_12_, per_din_13_, per_din_14_, per_din_15_, per_en, per_we_0_, per_we_1_, pmem_addr_0_, pmem_addr_1_, pmem_addr_2_, pmem_addr_3_, pmem_addr_4_, pmem_addr_5_, pmem_addr_6_, pmem_addr_7_, pmem_addr_8_, pmem_addr_9_, pmem_addr_10_, pmem_addr_11_, pmem_addr_12_, pmem_addr_13_, pmem_cen, pmem_din_0_, pmem_din_1_, pmem_din_2_, pmem_din_3_, pmem_din_4_, pmem_din_5_, pmem_din_6_, pmem_din_7_, pmem_din_8_, pmem_din_9_, pmem_din_10_, pmem_din_11_, pmem_din_12_, pmem_din_13_, pmem_din_14_, pmem_din_15_, pmem_wen_0_, pmem_wen_1_, puc_rst, smclk, smclk_en, cpu_en, dbg_en, dbg_i2c_addr_0_, dbg_i2c_addr_1_, dbg_i2c_addr_2_, dbg_i2c_addr_3_, dbg_i2c_addr_4_, dbg_i2c_addr_5_, dbg_i2c_addr_6_, dbg_i2c_broadcast_0_, dbg_i2c_broadcast_1_, dbg_i2c_broadcast_2_, dbg_i2c_broadcast_3_, dbg_i2c_broadcast_4_, dbg_i2c_broadcast_5_, dbg_i2c_broadcast_6_, dbg_i2c_scl, dbg_i2c_sda_in, dbg_uart_rxd, dco_clk, dmem_dout_0_, dmem_dout_1_, dmem_dout_2_, dmem_dout_3_, dmem_dout_4_, dmem_dout_5_, dmem_dout_6_, dmem_dout_7_, dmem_dout_8_, dmem_dout_9_, dmem_dout_10_, dmem_dout_11_, dmem_dout_12_, dmem_dout_13_, dmem_dout_14_, dmem_dout_15_, irq_0_, irq_1_, irq_2_, irq_3_, irq_4_, irq_5_, irq_6_, irq_7_, irq_8_, irq_9_, irq_10_, irq_11_, irq_12_, irq_13_, lfxt_clk, dma_addr_1_, dma_addr_2_, dma_addr_3_, dma_addr_4_, dma_addr_5_, dma_addr_6_, dma_addr_7_, dma_addr_8_, dma_addr_9_, dma_addr_10_, dma_addr_11_, dma_addr_12_, dma_addr_13_, dma_addr_14_, dma_addr_15_, dma_din_0_, dma_din_1_, dma_din_2_, dma_din_3_, dma_din_4_, dma_din_5_, dma_din_6_, dma_din_7_, dma_din_8_, dma_din_9_, dma_din_10_, dma_din_11_, dma_din_12_, dma_din_13_, dma_din_14_, dma_din_15_, dma_en, dma_priority, dma_we_0_, dma_we_1_, dma_wkup, nmi, per_dout_0_, per_dout_1_, per_dout_2_, per_dout_3_, per_dout_4_, per_dout_5_, per_dout_6_, per_dout_7_, per_dout_8_, per_dout_9_, per_dout_10_, per_dout_11_, per_dout_12_, per_dout_13_, per_dout_14_, per_dout_15_, pmem_dout_0_, pmem_dout_1_, pmem_dout_2_, pmem_dout_3_, pmem_dout_4_, pmem_dout_5_, pmem_dout_6_, pmem_dout_7_, pmem_dout_8_, pmem_dout_9_, pmem_dout_10_, pmem_dout_11_, pmem_dout_12_, pmem_dout_13_, pmem_dout_14_, pmem_dout_15_, reset_n, scan_enable, scan_mode, wkup);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire UNUSED_fe_mab_0;
  output aclk;
  output aclk_en;
  wire clock_module_0.UNUSED_cpuoff ;
  wire clock_module_0.aclk_div_0_ ;
  wire clock_module_0.aclk_div_1_ ;
  wire clock_module_0.aclk_div_2_ ;
  wire clock_module_0.bcsctl1_0_ ;
  wire clock_module_0.bcsctl1_1_ ;
  wire clock_module_0.bcsctl1_2_ ;
  wire clock_module_0.bcsctl1_3_ ;
  wire clock_module_0.bcsctl1_4_ ;
  wire clock_module_0.bcsctl1_5_ ;
  wire clock_module_0.bcsctl1_6_ ;
  wire clock_module_0.bcsctl1_7_ ;
  wire clock_module_0.bcsctl1_rd_10_ ;
  wire clock_module_0.bcsctl1_rd_11_ ;
  wire clock_module_0.bcsctl1_rd_12_ ;
  wire clock_module_0.bcsctl1_rd_13_ ;
  wire clock_module_0.bcsctl1_rd_14_ ;
  wire clock_module_0.bcsctl1_rd_15_ ;
  wire clock_module_0.bcsctl1_rd_8_ ;
  wire clock_module_0.bcsctl1_rd_9_ ;
  wire clock_module_0.bcsctl2_0_ ;
  wire clock_module_0.bcsctl2_1_ ;
  wire clock_module_0.bcsctl2_2_ ;
  wire clock_module_0.bcsctl2_3_ ;
  wire clock_module_0.bcsctl2_4_ ;
  wire clock_module_0.bcsctl2_5_ ;
  wire clock_module_0.bcsctl2_6_ ;
  wire clock_module_0.bcsctl2_7_ ;
  wire clock_module_0.bcsctl2_rd_0_ ;
  wire clock_module_0.bcsctl2_rd_1_ ;
  wire clock_module_0.bcsctl2_rd_2_ ;
  wire clock_module_0.bcsctl2_rd_3_ ;
  wire clock_module_0.bcsctl2_rd_4_ ;
  wire clock_module_0.bcsctl2_rd_5_ ;
  wire clock_module_0.bcsctl2_rd_6_ ;
  wire clock_module_0.bcsctl2_rd_7_ ;
  wire clock_module_0.dbg_cpu_reset ;
  wire clock_module_0.dbg_rst ;
  wire clock_module_0.dbg_rst_nxt ;
  wire clock_module_0.lfxt_clk_dly ;
  wire clock_module_0.lfxt_clk_s ;
  wire clock_module_0.oscoff ;
  wire clock_module_0.por ;
  wire clock_module_0.por_a ;
  wire clock_module_0.puc_a ;
  wire clock_module_0.puc_noscan_n ;
  wire clock_module_0.scg1 ;
  wire clock_module_0.smclk_div_0_ ;
  wire clock_module_0.smclk_div_1_ ;
  wire clock_module_0.smclk_div_2_ ;
  wire clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ;
  wire clock_module_0.sync_cell_puc.data_in ;
  wire clock_module_0.sync_cell_puc.data_sync_0_ ;
  wire clock_module_0.sync_reset_por.data_sync_0_ ;
  wire clock_module_0.wdt_reset ;
  input cpu_en;
  wire cpu_halt_cmd;
  wire cpu_halt_st;
  wire dbg_0.UNUSED_eu_mab_0_ ;
  wire dbg_0.UNUSED_eu_mab_10_ ;
  wire dbg_0.UNUSED_eu_mab_11_ ;
  wire dbg_0.UNUSED_eu_mab_12_ ;
  wire dbg_0.UNUSED_eu_mab_13_ ;
  wire dbg_0.UNUSED_eu_mab_14_ ;
  wire dbg_0.UNUSED_eu_mab_15_ ;
  wire dbg_0.UNUSED_eu_mab_1_ ;
  wire dbg_0.UNUSED_eu_mab_2_ ;
  wire dbg_0.UNUSED_eu_mab_3_ ;
  wire dbg_0.UNUSED_eu_mab_4_ ;
  wire dbg_0.UNUSED_eu_mab_5_ ;
  wire dbg_0.UNUSED_eu_mab_6_ ;
  wire dbg_0.UNUSED_eu_mab_7_ ;
  wire dbg_0.UNUSED_eu_mab_8_ ;
  wire dbg_0.UNUSED_eu_mab_9_ ;
  wire dbg_0.UNUSED_eu_mb_en ;
  wire dbg_0.UNUSED_eu_mb_wr_0_ ;
  wire dbg_0.UNUSED_eu_mb_wr_1_ ;
  wire dbg_0.UNUSED_pc_0_ ;
  wire dbg_0.UNUSED_pc_10_ ;
  wire dbg_0.UNUSED_pc_11_ ;
  wire dbg_0.UNUSED_pc_12_ ;
  wire dbg_0.UNUSED_pc_13_ ;
  wire dbg_0.UNUSED_pc_14_ ;
  wire dbg_0.UNUSED_pc_15_ ;
  wire dbg_0.UNUSED_pc_1_ ;
  wire dbg_0.UNUSED_pc_2_ ;
  wire dbg_0.UNUSED_pc_3_ ;
  wire dbg_0.UNUSED_pc_4_ ;
  wire dbg_0.UNUSED_pc_5_ ;
  wire dbg_0.UNUSED_pc_6_ ;
  wire dbg_0.UNUSED_pc_7_ ;
  wire dbg_0.UNUSED_pc_8_ ;
  wire dbg_0.UNUSED_pc_9_ ;
  wire dbg_0.cpu_ctl_3_ ;
  wire dbg_0.cpu_ctl_4_ ;
  wire dbg_0.cpu_ctl_5_ ;
  wire dbg_0.cpu_stat_2_ ;
  wire dbg_0.cpu_stat_3_ ;
  wire dbg_0.dbg_addr_0_ ;
  wire dbg_0.dbg_addr_1_ ;
  wire dbg_0.dbg_addr_2_ ;
  wire dbg_0.dbg_addr_3_ ;
  wire dbg_0.dbg_addr_4_ ;
  wire dbg_0.dbg_addr_5_ ;
  wire dbg_0.dbg_din_0_ ;
  wire dbg_0.dbg_din_10_ ;
  wire dbg_0.dbg_din_11_ ;
  wire dbg_0.dbg_din_12_ ;
  wire dbg_0.dbg_din_13_ ;
  wire dbg_0.dbg_din_14_ ;
  wire dbg_0.dbg_din_15_ ;
  wire dbg_0.dbg_din_1_ ;
  wire dbg_0.dbg_din_2_ ;
  wire dbg_0.dbg_din_3_ ;
  wire dbg_0.dbg_din_4_ ;
  wire dbg_0.dbg_din_5_ ;
  wire dbg_0.dbg_din_6_ ;
  wire dbg_0.dbg_din_7_ ;
  wire dbg_0.dbg_din_8_ ;
  wire dbg_0.dbg_din_9_ ;
  wire dbg_0.dbg_dout_0_ ;
  wire dbg_0.dbg_dout_10_ ;
  wire dbg_0.dbg_dout_11_ ;
  wire dbg_0.dbg_dout_12_ ;
  wire dbg_0.dbg_dout_13_ ;
  wire dbg_0.dbg_dout_14_ ;
  wire dbg_0.dbg_dout_15_ ;
  wire dbg_0.dbg_dout_1_ ;
  wire dbg_0.dbg_dout_2_ ;
  wire dbg_0.dbg_dout_3_ ;
  wire dbg_0.dbg_dout_4_ ;
  wire dbg_0.dbg_dout_5_ ;
  wire dbg_0.dbg_dout_6_ ;
  wire dbg_0.dbg_dout_7_ ;
  wire dbg_0.dbg_dout_8_ ;
  wire dbg_0.dbg_dout_9_ ;
  wire dbg_0.dbg_i2c_0.dbg_bw ;
  wire dbg_0.dbg_i2c_0.dbg_rd ;
  wire dbg_0.dbg_i2c_0.dbg_state_0_ ;
  wire dbg_0.dbg_i2c_0.dbg_state_1_ ;
  wire dbg_0.dbg_i2c_0.dbg_state_2_ ;
  wire dbg_0.dbg_i2c_0.dbg_state_3_ ;
  wire dbg_0.dbg_i2c_0.dbg_state_4_ ;
  wire dbg_0.dbg_i2c_0.dbg_wr ;
  wire dbg_0.dbg_i2c_0.i2c_active_seq ;
  wire dbg_0.dbg_i2c_0.i2c_state_0_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_1_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_2_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_3_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_4_ ;
  wire dbg_0.dbg_i2c_0.i2c_state_5_ ;
  wire dbg_0.dbg_i2c_0.mem_burst ;
  wire dbg_0.dbg_i2c_0.mem_burst_end ;
  wire dbg_0.dbg_i2c_0.mem_burst_rd ;
  wire dbg_0.dbg_i2c_0.mem_burst_wr ;
  wire dbg_0.dbg_i2c_0.mem_bw ;
  wire dbg_0.dbg_i2c_0.scl ;
  wire dbg_0.dbg_i2c_0.scl_buf_0_ ;
  wire dbg_0.dbg_i2c_0.scl_buf_1_ ;
  wire dbg_0.dbg_i2c_0.scl_dly ;
  wire dbg_0.dbg_i2c_0.scl_re ;
  wire dbg_0.dbg_i2c_0.scl_re_dly_0_ ;
  wire dbg_0.dbg_i2c_0.scl_re_dly_1_ ;
  wire dbg_0.dbg_i2c_0.scl_sync ;
  wire dbg_0.dbg_i2c_0.scl_sync_n ;
  wire dbg_0.dbg_i2c_0.sda_in ;
  wire dbg_0.dbg_i2c_0.sda_in_buf_0_ ;
  wire dbg_0.dbg_i2c_0.sda_in_buf_1_ ;
  wire dbg_0.dbg_i2c_0.sda_in_dly ;
  wire dbg_0.dbg_i2c_0.sda_in_sync ;
  wire dbg_0.dbg_i2c_0.sda_in_sync_n ;
  wire dbg_0.dbg_i2c_0.shift_buf_0_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_1_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_2_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_3_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_4_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_5_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_6_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_7_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_8_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_0_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_1_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_2_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_3_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_4_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_5_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_6_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_7_ ;
  wire dbg_0.dbg_i2c_0.shift_buf_nxt_8_ ;
  wire dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in ;
  wire dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ;
  wire dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in ;
  wire dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ;
  wire dbg_0.dbg_mem_addr_0_ ;
  wire dbg_0.dbg_mem_addr_10_ ;
  wire dbg_0.dbg_mem_addr_11_ ;
  wire dbg_0.dbg_mem_addr_12_ ;
  wire dbg_0.dbg_mem_addr_13_ ;
  wire dbg_0.dbg_mem_addr_14_ ;
  wire dbg_0.dbg_mem_addr_15_ ;
  wire dbg_0.dbg_mem_addr_1_ ;
  wire dbg_0.dbg_mem_addr_2_ ;
  wire dbg_0.dbg_mem_addr_3_ ;
  wire dbg_0.dbg_mem_addr_4_ ;
  wire dbg_0.dbg_mem_addr_5_ ;
  wire dbg_0.dbg_mem_addr_6_ ;
  wire dbg_0.dbg_mem_addr_7_ ;
  wire dbg_0.dbg_mem_addr_8_ ;
  wire dbg_0.dbg_mem_addr_9_ ;
  wire dbg_0.dbg_mem_din_0_ ;
  wire dbg_0.dbg_mem_din_10_ ;
  wire dbg_0.dbg_mem_din_11_ ;
  wire dbg_0.dbg_mem_din_12_ ;
  wire dbg_0.dbg_mem_din_13_ ;
  wire dbg_0.dbg_mem_din_14_ ;
  wire dbg_0.dbg_mem_din_15_ ;
  wire dbg_0.dbg_mem_din_1_ ;
  wire dbg_0.dbg_mem_din_2_ ;
  wire dbg_0.dbg_mem_din_3_ ;
  wire dbg_0.dbg_mem_din_4_ ;
  wire dbg_0.dbg_mem_din_5_ ;
  wire dbg_0.dbg_mem_din_6_ ;
  wire dbg_0.dbg_mem_din_7_ ;
  wire dbg_0.dbg_mem_din_8_ ;
  wire dbg_0.dbg_mem_din_9_ ;
  wire dbg_0.dbg_mem_en ;
  wire dbg_0.dbg_mem_rd ;
  wire dbg_0.dbg_mem_rd_dly ;
  wire dbg_0.dbg_mem_wr_0_ ;
  wire dbg_0.dbg_mem_wr_1_ ;
  wire dbg_0.dbg_rd_rdy ;
  wire dbg_0.dbg_reg_din_0_ ;
  wire dbg_0.dbg_reg_din_10_ ;
  wire dbg_0.dbg_reg_din_11_ ;
  wire dbg_0.dbg_reg_din_12_ ;
  wire dbg_0.dbg_reg_din_13_ ;
  wire dbg_0.dbg_reg_din_14_ ;
  wire dbg_0.dbg_reg_din_15_ ;
  wire dbg_0.dbg_reg_din_1_ ;
  wire dbg_0.dbg_reg_din_2_ ;
  wire dbg_0.dbg_reg_din_3_ ;
  wire dbg_0.dbg_reg_din_4_ ;
  wire dbg_0.dbg_reg_din_5_ ;
  wire dbg_0.dbg_reg_din_6_ ;
  wire dbg_0.dbg_reg_din_7_ ;
  wire dbg_0.dbg_reg_din_8_ ;
  wire dbg_0.dbg_reg_din_9_ ;
  wire dbg_0.dbg_reg_wr ;
  wire dbg_0.decode_noirq ;
  wire dbg_0.fe_mdb_in_0_ ;
  wire dbg_0.fe_mdb_in_10_ ;
  wire dbg_0.fe_mdb_in_11_ ;
  wire dbg_0.fe_mdb_in_12_ ;
  wire dbg_0.fe_mdb_in_13_ ;
  wire dbg_0.fe_mdb_in_14_ ;
  wire dbg_0.fe_mdb_in_15_ ;
  wire dbg_0.fe_mdb_in_1_ ;
  wire dbg_0.fe_mdb_in_2_ ;
  wire dbg_0.fe_mdb_in_3_ ;
  wire dbg_0.fe_mdb_in_4_ ;
  wire dbg_0.fe_mdb_in_5_ ;
  wire dbg_0.fe_mdb_in_6_ ;
  wire dbg_0.fe_mdb_in_7_ ;
  wire dbg_0.fe_mdb_in_8_ ;
  wire dbg_0.fe_mdb_in_9_ ;
  wire dbg_0.halt_flag ;
  wire dbg_0.inc_step_0_ ;
  wire dbg_0.inc_step_1_ ;
  wire dbg_0.istep ;
  wire dbg_0.mem_cnt_0_ ;
  wire dbg_0.mem_cnt_10_ ;
  wire dbg_0.mem_cnt_11_ ;
  wire dbg_0.mem_cnt_12_ ;
  wire dbg_0.mem_cnt_13_ ;
  wire dbg_0.mem_cnt_14_ ;
  wire dbg_0.mem_cnt_15_ ;
  wire dbg_0.mem_cnt_1_ ;
  wire dbg_0.mem_cnt_2_ ;
  wire dbg_0.mem_cnt_3_ ;
  wire dbg_0.mem_cnt_4_ ;
  wire dbg_0.mem_cnt_5_ ;
  wire dbg_0.mem_cnt_6_ ;
  wire dbg_0.mem_cnt_7_ ;
  wire dbg_0.mem_cnt_8_ ;
  wire dbg_0.mem_cnt_9_ ;
  wire dbg_0.mem_ctl_1_ ;
  wire dbg_0.mem_ctl_2_ ;
  wire dbg_0.mem_data_0_ ;
  wire dbg_0.mem_data_10_ ;
  wire dbg_0.mem_data_11_ ;
  wire dbg_0.mem_data_12_ ;
  wire dbg_0.mem_data_13_ ;
  wire dbg_0.mem_data_14_ ;
  wire dbg_0.mem_data_15_ ;
  wire dbg_0.mem_data_1_ ;
  wire dbg_0.mem_data_2_ ;
  wire dbg_0.mem_data_3_ ;
  wire dbg_0.mem_data_4_ ;
  wire dbg_0.mem_data_5_ ;
  wire dbg_0.mem_data_6_ ;
  wire dbg_0.mem_data_7_ ;
  wire dbg_0.mem_data_8_ ;
  wire dbg_0.mem_data_9_ ;
  wire dbg_0.mem_start ;
  wire dbg_0.mem_startb ;
  wire dbg_0.mem_state_0_ ;
  wire dbg_0.mem_state_1_ ;
  wire dbg_0.mem_state_2_ ;
  wire dbg_0.mem_state_3_ ;
  input dbg_en;
  output dbg_freeze;
  input dbg_i2c_addr_0_;
  input dbg_i2c_addr_1_;
  input dbg_i2c_addr_2_;
  input dbg_i2c_addr_3_;
  input dbg_i2c_addr_4_;
  input dbg_i2c_addr_5_;
  input dbg_i2c_addr_6_;
  input dbg_i2c_broadcast_0_;
  input dbg_i2c_broadcast_1_;
  input dbg_i2c_broadcast_2_;
  input dbg_i2c_broadcast_3_;
  input dbg_i2c_broadcast_4_;
  input dbg_i2c_broadcast_5_;
  input dbg_i2c_broadcast_6_;
  input dbg_i2c_scl;
  input dbg_i2c_sda_in;
  output dbg_i2c_sda_out;
  input dbg_uart_rxd;
  output dbg_uart_txd;
  input dco_clk;
  output dco_enable;
  output dco_wkup;
  input dma_addr_10_;
  input dma_addr_11_;
  input dma_addr_12_;
  input dma_addr_13_;
  input dma_addr_14_;
  input dma_addr_15_;
  input dma_addr_1_;
  input dma_addr_2_;
  input dma_addr_3_;
  input dma_addr_4_;
  input dma_addr_5_;
  input dma_addr_6_;
  input dma_addr_7_;
  input dma_addr_8_;
  input dma_addr_9_;
  input dma_din_0_;
  input dma_din_10_;
  input dma_din_11_;
  input dma_din_12_;
  input dma_din_13_;
  input dma_din_14_;
  input dma_din_15_;
  input dma_din_1_;
  input dma_din_2_;
  input dma_din_3_;
  input dma_din_4_;
  input dma_din_5_;
  input dma_din_6_;
  input dma_din_7_;
  input dma_din_8_;
  input dma_din_9_;
  output dma_dout_0_;
  output dma_dout_10_;
  output dma_dout_11_;
  output dma_dout_12_;
  output dma_dout_13_;
  output dma_dout_14_;
  output dma_dout_15_;
  output dma_dout_1_;
  output dma_dout_2_;
  output dma_dout_3_;
  output dma_dout_4_;
  output dma_dout_5_;
  output dma_dout_6_;
  output dma_dout_7_;
  output dma_dout_8_;
  output dma_dout_9_;
  input dma_en;
  input dma_priority;
  output dma_ready;
  output dma_resp;
  input dma_we_0_;
  input dma_we_1_;
  input dma_wkup;
  output dmem_addr_0_;
  output dmem_addr_10_;
  output dmem_addr_11_;
  output dmem_addr_12_;
  output dmem_addr_1_;
  output dmem_addr_2_;
  output dmem_addr_3_;
  output dmem_addr_4_;
  output dmem_addr_5_;
  output dmem_addr_6_;
  output dmem_addr_7_;
  output dmem_addr_8_;
  output dmem_addr_9_;
  output dmem_cen;
  output dmem_din_0_;
  output dmem_din_10_;
  output dmem_din_11_;
  output dmem_din_12_;
  output dmem_din_13_;
  output dmem_din_14_;
  output dmem_din_15_;
  output dmem_din_1_;
  output dmem_din_2_;
  output dmem_din_3_;
  output dmem_din_4_;
  output dmem_din_5_;
  output dmem_din_6_;
  output dmem_din_7_;
  output dmem_din_8_;
  output dmem_din_9_;
  input dmem_dout_0_;
  input dmem_dout_10_;
  input dmem_dout_11_;
  input dmem_dout_12_;
  input dmem_dout_13_;
  input dmem_dout_14_;
  input dmem_dout_15_;
  input dmem_dout_1_;
  input dmem_dout_2_;
  input dmem_dout_3_;
  input dmem_dout_4_;
  input dmem_dout_5_;
  input dmem_dout_6_;
  input dmem_dout_7_;
  input dmem_dout_8_;
  input dmem_dout_9_;
  output dmem_wen_0_;
  output dmem_wen_1_;
  wire e_state_0_;
  wire e_state_1_;
  wire e_state_2_;
  wire e_state_3_;
  wire eu_mdb_in_0_;
  wire eu_mdb_in_10_;
  wire eu_mdb_in_11_;
  wire eu_mdb_in_12_;
  wire eu_mdb_in_13_;
  wire eu_mdb_in_14_;
  wire eu_mdb_in_15_;
  wire eu_mdb_in_1_;
  wire eu_mdb_in_2_;
  wire eu_mdb_in_3_;
  wire eu_mdb_in_4_;
  wire eu_mdb_in_5_;
  wire eu_mdb_in_6_;
  wire eu_mdb_in_7_;
  wire eu_mdb_in_8_;
  wire eu_mdb_in_9_;
  wire eu_mdb_out_0_;
  wire eu_mdb_out_10_;
  wire eu_mdb_out_11_;
  wire eu_mdb_out_12_;
  wire eu_mdb_out_13_;
  wire eu_mdb_out_14_;
  wire eu_mdb_out_15_;
  wire eu_mdb_out_1_;
  wire eu_mdb_out_2_;
  wire eu_mdb_out_3_;
  wire eu_mdb_out_4_;
  wire eu_mdb_out_5_;
  wire eu_mdb_out_6_;
  wire eu_mdb_out_7_;
  wire eu_mdb_out_8_;
  wire eu_mdb_out_9_;
  wire exec_done;
  wire execution_unit_0.UNUSED_inst_ad_idx ;
  wire execution_unit_0.UNUSED_inst_ad_symb ;
  wire execution_unit_0.alu_0.N ;
  wire execution_unit_0.alu_0.UNUSED_inst_alu ;
  wire execution_unit_0.alu_0.UNUSED_inst_so_call ;
  wire execution_unit_0.alu_0.UNUSED_inst_so_push ;
  wire execution_unit_0.alu_0.UNUSED_inst_so_reti ;
  wire execution_unit_0.alu_0.Z ;
  wire execution_unit_0.alu_0.alu_out_0_ ;
  wire execution_unit_0.alu_0.alu_out_10_ ;
  wire execution_unit_0.alu_0.alu_out_11_ ;
  wire execution_unit_0.alu_0.alu_out_12_ ;
  wire execution_unit_0.alu_0.alu_out_13_ ;
  wire execution_unit_0.alu_0.alu_out_14_ ;
  wire execution_unit_0.alu_0.alu_out_15_ ;
  wire execution_unit_0.alu_0.alu_out_1_ ;
  wire execution_unit_0.alu_0.alu_out_2_ ;
  wire execution_unit_0.alu_0.alu_out_3_ ;
  wire execution_unit_0.alu_0.alu_out_4_ ;
  wire execution_unit_0.alu_0.alu_out_5_ ;
  wire execution_unit_0.alu_0.alu_out_6_ ;
  wire execution_unit_0.alu_0.alu_out_7_ ;
  wire execution_unit_0.alu_0.alu_out_8_ ;
  wire execution_unit_0.alu_0.alu_out_9_ ;
  wire execution_unit_0.alu_0.alu_shift_0_ ;
  wire execution_unit_0.alu_0.alu_shift_10_ ;
  wire execution_unit_0.alu_0.alu_shift_11_ ;
  wire execution_unit_0.alu_0.alu_shift_12_ ;
  wire execution_unit_0.alu_0.alu_shift_13_ ;
  wire execution_unit_0.alu_0.alu_shift_14_ ;
  wire execution_unit_0.alu_0.alu_shift_1_ ;
  wire execution_unit_0.alu_0.alu_shift_2_ ;
  wire execution_unit_0.alu_0.alu_shift_3_ ;
  wire execution_unit_0.alu_0.alu_shift_4_ ;
  wire execution_unit_0.alu_0.alu_shift_5_ ;
  wire execution_unit_0.alu_0.alu_shift_6_ ;
  wire execution_unit_0.alu_0.alu_shift_8_ ;
  wire execution_unit_0.alu_0.alu_shift_9_ ;
  wire execution_unit_0.alu_0.alu_stat_0_ ;
  wire execution_unit_0.alu_0.alu_stat_3_ ;
  wire execution_unit_0.alu_0.alu_stat_wr_0_ ;
  wire execution_unit_0.alu_0.alu_swpb_0_ ;
  wire execution_unit_0.alu_0.alu_swpb_8_ ;
  wire execution_unit_0.alu_0.exec_cycle ;
  wire execution_unit_0.alu_0.inst_alu_0_ ;
  wire execution_unit_0.alu_0.inst_alu_10_ ;
  wire execution_unit_0.alu_0.inst_alu_1_ ;
  wire execution_unit_0.alu_0.inst_alu_2_ ;
  wire execution_unit_0.alu_0.inst_alu_3_ ;
  wire execution_unit_0.alu_0.inst_alu_4_ ;
  wire execution_unit_0.alu_0.inst_alu_5_ ;
  wire execution_unit_0.alu_0.inst_alu_6_ ;
  wire execution_unit_0.alu_0.inst_alu_7_ ;
  wire execution_unit_0.alu_0.inst_alu_8_ ;
  wire execution_unit_0.alu_0.inst_alu_9_ ;
  wire execution_unit_0.alu_0.inst_bw ;
  wire execution_unit_0.alu_0.inst_jmp_0_ ;
  wire execution_unit_0.alu_0.inst_jmp_1_ ;
  wire execution_unit_0.alu_0.inst_jmp_2_ ;
  wire execution_unit_0.alu_0.inst_jmp_3_ ;
  wire execution_unit_0.alu_0.inst_jmp_4_ ;
  wire execution_unit_0.alu_0.inst_jmp_5_ ;
  wire execution_unit_0.alu_0.inst_jmp_6_ ;
  wire execution_unit_0.alu_0.inst_so_0_ ;
  wire execution_unit_0.alu_0.inst_so_1_ ;
  wire execution_unit_0.alu_0.inst_so_3_ ;
  wire execution_unit_0.alu_0.inst_so_7_ ;
  wire execution_unit_0.alu_0.op_dst_0_ ;
  wire execution_unit_0.alu_0.op_dst_10_ ;
  wire execution_unit_0.alu_0.op_dst_11_ ;
  wire execution_unit_0.alu_0.op_dst_12_ ;
  wire execution_unit_0.alu_0.op_dst_13_ ;
  wire execution_unit_0.alu_0.op_dst_14_ ;
  wire execution_unit_0.alu_0.op_dst_15_ ;
  wire execution_unit_0.alu_0.op_dst_1_ ;
  wire execution_unit_0.alu_0.op_dst_2_ ;
  wire execution_unit_0.alu_0.op_dst_3_ ;
  wire execution_unit_0.alu_0.op_dst_4_ ;
  wire execution_unit_0.alu_0.op_dst_5_ ;
  wire execution_unit_0.alu_0.op_dst_6_ ;
  wire execution_unit_0.alu_0.op_dst_7_ ;
  wire execution_unit_0.alu_0.op_dst_8_ ;
  wire execution_unit_0.alu_0.op_dst_9_ ;
  wire execution_unit_0.alu_0.status_0_ ;
  wire execution_unit_0.alu_0.status_1_ ;
  wire execution_unit_0.alu_0.status_2_ ;
  wire execution_unit_0.alu_0.status_3_ ;
  wire execution_unit_0.gie ;
  wire execution_unit_0.inst_ad_0_ ;
  wire execution_unit_0.inst_ad_6_ ;
  wire execution_unit_0.inst_as_0_ ;
  wire execution_unit_0.inst_as_1_ ;
  wire execution_unit_0.inst_as_2_ ;
  wire execution_unit_0.inst_as_3_ ;
  wire execution_unit_0.inst_as_4_ ;
  wire execution_unit_0.inst_as_5_ ;
  wire execution_unit_0.inst_as_6_ ;
  wire execution_unit_0.inst_as_7_ ;
  wire execution_unit_0.inst_dest_0_ ;
  wire execution_unit_0.inst_dest_10_ ;
  wire execution_unit_0.inst_dest_11_ ;
  wire execution_unit_0.inst_dest_12_ ;
  wire execution_unit_0.inst_dest_13_ ;
  wire execution_unit_0.inst_dest_14_ ;
  wire execution_unit_0.inst_dest_15_ ;
  wire execution_unit_0.inst_dest_1_ ;
  wire execution_unit_0.inst_dest_2_ ;
  wire execution_unit_0.inst_dest_3_ ;
  wire execution_unit_0.inst_dest_4_ ;
  wire execution_unit_0.inst_dest_5_ ;
  wire execution_unit_0.inst_dest_6_ ;
  wire execution_unit_0.inst_dest_7_ ;
  wire execution_unit_0.inst_dest_8_ ;
  wire execution_unit_0.inst_dest_9_ ;
  wire execution_unit_0.inst_dext_0_ ;
  wire execution_unit_0.inst_dext_10_ ;
  wire execution_unit_0.inst_dext_11_ ;
  wire execution_unit_0.inst_dext_12_ ;
  wire execution_unit_0.inst_dext_13_ ;
  wire execution_unit_0.inst_dext_14_ ;
  wire execution_unit_0.inst_dext_15_ ;
  wire execution_unit_0.inst_dext_1_ ;
  wire execution_unit_0.inst_dext_2_ ;
  wire execution_unit_0.inst_dext_3_ ;
  wire execution_unit_0.inst_dext_4_ ;
  wire execution_unit_0.inst_dext_5_ ;
  wire execution_unit_0.inst_dext_6_ ;
  wire execution_unit_0.inst_dext_7_ ;
  wire execution_unit_0.inst_dext_8_ ;
  wire execution_unit_0.inst_dext_9_ ;
  wire execution_unit_0.inst_irq_rst ;
  wire execution_unit_0.inst_mov ;
  wire execution_unit_0.inst_sext_0_ ;
  wire execution_unit_0.inst_sext_10_ ;
  wire execution_unit_0.inst_sext_11_ ;
  wire execution_unit_0.inst_sext_12_ ;
  wire execution_unit_0.inst_sext_13_ ;
  wire execution_unit_0.inst_sext_14_ ;
  wire execution_unit_0.inst_sext_15_ ;
  wire execution_unit_0.inst_sext_1_ ;
  wire execution_unit_0.inst_sext_2_ ;
  wire execution_unit_0.inst_sext_3_ ;
  wire execution_unit_0.inst_sext_4_ ;
  wire execution_unit_0.inst_sext_5_ ;
  wire execution_unit_0.inst_sext_6_ ;
  wire execution_unit_0.inst_sext_7_ ;
  wire execution_unit_0.inst_sext_8_ ;
  wire execution_unit_0.inst_sext_9_ ;
  wire execution_unit_0.inst_src_0_ ;
  wire execution_unit_0.inst_src_10_ ;
  wire execution_unit_0.inst_src_11_ ;
  wire execution_unit_0.inst_src_12_ ;
  wire execution_unit_0.inst_src_13_ ;
  wire execution_unit_0.inst_src_14_ ;
  wire execution_unit_0.inst_src_15_ ;
  wire execution_unit_0.inst_src_1_ ;
  wire execution_unit_0.inst_src_2_ ;
  wire execution_unit_0.inst_src_3_ ;
  wire execution_unit_0.inst_src_4_ ;
  wire execution_unit_0.inst_src_5_ ;
  wire execution_unit_0.inst_src_6_ ;
  wire execution_unit_0.inst_src_7_ ;
  wire execution_unit_0.inst_src_8_ ;
  wire execution_unit_0.inst_src_9_ ;
  wire execution_unit_0.inst_type_0_ ;
  wire execution_unit_0.inst_type_1_ ;
  wire execution_unit_0.inst_type_2_ ;
  wire execution_unit_0.mab_lsb ;
  wire execution_unit_0.mdb_in_buf_0_ ;
  wire execution_unit_0.mdb_in_buf_10_ ;
  wire execution_unit_0.mdb_in_buf_11_ ;
  wire execution_unit_0.mdb_in_buf_12_ ;
  wire execution_unit_0.mdb_in_buf_13_ ;
  wire execution_unit_0.mdb_in_buf_14_ ;
  wire execution_unit_0.mdb_in_buf_15_ ;
  wire execution_unit_0.mdb_in_buf_1_ ;
  wire execution_unit_0.mdb_in_buf_2_ ;
  wire execution_unit_0.mdb_in_buf_3_ ;
  wire execution_unit_0.mdb_in_buf_4_ ;
  wire execution_unit_0.mdb_in_buf_5_ ;
  wire execution_unit_0.mdb_in_buf_6_ ;
  wire execution_unit_0.mdb_in_buf_7_ ;
  wire execution_unit_0.mdb_in_buf_8_ ;
  wire execution_unit_0.mdb_in_buf_9_ ;
  wire execution_unit_0.mdb_in_buf_en ;
  wire execution_unit_0.mdb_in_buf_valid ;
  wire execution_unit_0.mdb_out_nxt_10_ ;
  wire execution_unit_0.mdb_out_nxt_11_ ;
  wire execution_unit_0.mdb_out_nxt_12_ ;
  wire execution_unit_0.mdb_out_nxt_13_ ;
  wire execution_unit_0.mdb_out_nxt_14_ ;
  wire execution_unit_0.mdb_out_nxt_15_ ;
  wire execution_unit_0.mdb_out_nxt_8_ ;
  wire execution_unit_0.mdb_out_nxt_9_ ;
  wire execution_unit_0.pc_nxt_10_ ;
  wire execution_unit_0.pc_nxt_11_ ;
  wire execution_unit_0.pc_nxt_12_ ;
  wire execution_unit_0.pc_nxt_13_ ;
  wire execution_unit_0.pc_nxt_14_ ;
  wire execution_unit_0.pc_nxt_15_ ;
  wire execution_unit_0.pc_nxt_1_ ;
  wire execution_unit_0.pc_nxt_2_ ;
  wire execution_unit_0.pc_nxt_3_ ;
  wire execution_unit_0.pc_nxt_4_ ;
  wire execution_unit_0.pc_nxt_5_ ;
  wire execution_unit_0.pc_nxt_6_ ;
  wire execution_unit_0.pc_nxt_7_ ;
  wire execution_unit_0.pc_nxt_8_ ;
  wire execution_unit_0.pc_nxt_9_ ;
  wire execution_unit_0.pc_sw_10_ ;
  wire execution_unit_0.pc_sw_11_ ;
  wire execution_unit_0.pc_sw_12_ ;
  wire execution_unit_0.pc_sw_13_ ;
  wire execution_unit_0.pc_sw_14_ ;
  wire execution_unit_0.pc_sw_15_ ;
  wire execution_unit_0.pc_sw_8_ ;
  wire execution_unit_0.pc_sw_9_ ;
  wire execution_unit_0.pc_sw_wr ;
  wire execution_unit_0.reg_dest_wr ;
  wire execution_unit_0.reg_incr ;
  wire execution_unit_0.reg_pc_call ;
  wire execution_unit_0.reg_sp_wr ;
  wire execution_unit_0.reg_sr_clr ;
  wire execution_unit_0.reg_sr_wr ;
  wire execution_unit_0.reg_src_0_ ;
  wire execution_unit_0.reg_src_10_ ;
  wire execution_unit_0.reg_src_11_ ;
  wire execution_unit_0.reg_src_12_ ;
  wire execution_unit_0.reg_src_13_ ;
  wire execution_unit_0.reg_src_14_ ;
  wire execution_unit_0.reg_src_15_ ;
  wire execution_unit_0.reg_src_1_ ;
  wire execution_unit_0.reg_src_2_ ;
  wire execution_unit_0.reg_src_3_ ;
  wire execution_unit_0.reg_src_4_ ;
  wire execution_unit_0.reg_src_5_ ;
  wire execution_unit_0.reg_src_6_ ;
  wire execution_unit_0.reg_src_7_ ;
  wire execution_unit_0.reg_src_8_ ;
  wire execution_unit_0.reg_src_9_ ;
  wire execution_unit_0.register_file_0.r10_0_ ;
  wire execution_unit_0.register_file_0.r10_10_ ;
  wire execution_unit_0.register_file_0.r10_11_ ;
  wire execution_unit_0.register_file_0.r10_12_ ;
  wire execution_unit_0.register_file_0.r10_13_ ;
  wire execution_unit_0.register_file_0.r10_14_ ;
  wire execution_unit_0.register_file_0.r10_15_ ;
  wire execution_unit_0.register_file_0.r10_1_ ;
  wire execution_unit_0.register_file_0.r10_2_ ;
  wire execution_unit_0.register_file_0.r10_3_ ;
  wire execution_unit_0.register_file_0.r10_4_ ;
  wire execution_unit_0.register_file_0.r10_5_ ;
  wire execution_unit_0.register_file_0.r10_6_ ;
  wire execution_unit_0.register_file_0.r10_7_ ;
  wire execution_unit_0.register_file_0.r10_8_ ;
  wire execution_unit_0.register_file_0.r10_9_ ;
  wire execution_unit_0.register_file_0.r11_0_ ;
  wire execution_unit_0.register_file_0.r11_10_ ;
  wire execution_unit_0.register_file_0.r11_11_ ;
  wire execution_unit_0.register_file_0.r11_12_ ;
  wire execution_unit_0.register_file_0.r11_13_ ;
  wire execution_unit_0.register_file_0.r11_14_ ;
  wire execution_unit_0.register_file_0.r11_15_ ;
  wire execution_unit_0.register_file_0.r11_1_ ;
  wire execution_unit_0.register_file_0.r11_2_ ;
  wire execution_unit_0.register_file_0.r11_3_ ;
  wire execution_unit_0.register_file_0.r11_4_ ;
  wire execution_unit_0.register_file_0.r11_5_ ;
  wire execution_unit_0.register_file_0.r11_6_ ;
  wire execution_unit_0.register_file_0.r11_7_ ;
  wire execution_unit_0.register_file_0.r11_8_ ;
  wire execution_unit_0.register_file_0.r11_9_ ;
  wire execution_unit_0.register_file_0.r12_0_ ;
  wire execution_unit_0.register_file_0.r12_10_ ;
  wire execution_unit_0.register_file_0.r12_11_ ;
  wire execution_unit_0.register_file_0.r12_12_ ;
  wire execution_unit_0.register_file_0.r12_13_ ;
  wire execution_unit_0.register_file_0.r12_14_ ;
  wire execution_unit_0.register_file_0.r12_15_ ;
  wire execution_unit_0.register_file_0.r12_1_ ;
  wire execution_unit_0.register_file_0.r12_2_ ;
  wire execution_unit_0.register_file_0.r12_3_ ;
  wire execution_unit_0.register_file_0.r12_4_ ;
  wire execution_unit_0.register_file_0.r12_5_ ;
  wire execution_unit_0.register_file_0.r12_6_ ;
  wire execution_unit_0.register_file_0.r12_7_ ;
  wire execution_unit_0.register_file_0.r12_8_ ;
  wire execution_unit_0.register_file_0.r12_9_ ;
  wire execution_unit_0.register_file_0.r13_0_ ;
  wire execution_unit_0.register_file_0.r13_10_ ;
  wire execution_unit_0.register_file_0.r13_11_ ;
  wire execution_unit_0.register_file_0.r13_12_ ;
  wire execution_unit_0.register_file_0.r13_13_ ;
  wire execution_unit_0.register_file_0.r13_14_ ;
  wire execution_unit_0.register_file_0.r13_15_ ;
  wire execution_unit_0.register_file_0.r13_1_ ;
  wire execution_unit_0.register_file_0.r13_2_ ;
  wire execution_unit_0.register_file_0.r13_3_ ;
  wire execution_unit_0.register_file_0.r13_4_ ;
  wire execution_unit_0.register_file_0.r13_5_ ;
  wire execution_unit_0.register_file_0.r13_6_ ;
  wire execution_unit_0.register_file_0.r13_7_ ;
  wire execution_unit_0.register_file_0.r13_8_ ;
  wire execution_unit_0.register_file_0.r13_9_ ;
  wire execution_unit_0.register_file_0.r14_0_ ;
  wire execution_unit_0.register_file_0.r14_10_ ;
  wire execution_unit_0.register_file_0.r14_11_ ;
  wire execution_unit_0.register_file_0.r14_12_ ;
  wire execution_unit_0.register_file_0.r14_13_ ;
  wire execution_unit_0.register_file_0.r14_14_ ;
  wire execution_unit_0.register_file_0.r14_15_ ;
  wire execution_unit_0.register_file_0.r14_1_ ;
  wire execution_unit_0.register_file_0.r14_2_ ;
  wire execution_unit_0.register_file_0.r14_3_ ;
  wire execution_unit_0.register_file_0.r14_4_ ;
  wire execution_unit_0.register_file_0.r14_5_ ;
  wire execution_unit_0.register_file_0.r14_6_ ;
  wire execution_unit_0.register_file_0.r14_7_ ;
  wire execution_unit_0.register_file_0.r14_8_ ;
  wire execution_unit_0.register_file_0.r14_9_ ;
  wire execution_unit_0.register_file_0.r15_0_ ;
  wire execution_unit_0.register_file_0.r15_10_ ;
  wire execution_unit_0.register_file_0.r15_11_ ;
  wire execution_unit_0.register_file_0.r15_12_ ;
  wire execution_unit_0.register_file_0.r15_13_ ;
  wire execution_unit_0.register_file_0.r15_14_ ;
  wire execution_unit_0.register_file_0.r15_15_ ;
  wire execution_unit_0.register_file_0.r15_1_ ;
  wire execution_unit_0.register_file_0.r15_2_ ;
  wire execution_unit_0.register_file_0.r15_3_ ;
  wire execution_unit_0.register_file_0.r15_4_ ;
  wire execution_unit_0.register_file_0.r15_5_ ;
  wire execution_unit_0.register_file_0.r15_6_ ;
  wire execution_unit_0.register_file_0.r15_7_ ;
  wire execution_unit_0.register_file_0.r15_8_ ;
  wire execution_unit_0.register_file_0.r15_9_ ;
  wire execution_unit_0.register_file_0.r1_0_ ;
  wire execution_unit_0.register_file_0.r1_10_ ;
  wire execution_unit_0.register_file_0.r1_11_ ;
  wire execution_unit_0.register_file_0.r1_12_ ;
  wire execution_unit_0.register_file_0.r1_13_ ;
  wire execution_unit_0.register_file_0.r1_14_ ;
  wire execution_unit_0.register_file_0.r1_15_ ;
  wire execution_unit_0.register_file_0.r1_1_ ;
  wire execution_unit_0.register_file_0.r1_2_ ;
  wire execution_unit_0.register_file_0.r1_3_ ;
  wire execution_unit_0.register_file_0.r1_4_ ;
  wire execution_unit_0.register_file_0.r1_5_ ;
  wire execution_unit_0.register_file_0.r1_6_ ;
  wire execution_unit_0.register_file_0.r1_7_ ;
  wire execution_unit_0.register_file_0.r1_8_ ;
  wire execution_unit_0.register_file_0.r1_9_ ;
  wire execution_unit_0.register_file_0.r2_4_ ;
  wire execution_unit_0.register_file_0.r3_0_ ;
  wire execution_unit_0.register_file_0.r3_10_ ;
  wire execution_unit_0.register_file_0.r3_11_ ;
  wire execution_unit_0.register_file_0.r3_12_ ;
  wire execution_unit_0.register_file_0.r3_13_ ;
  wire execution_unit_0.register_file_0.r3_14_ ;
  wire execution_unit_0.register_file_0.r3_15_ ;
  wire execution_unit_0.register_file_0.r3_1_ ;
  wire execution_unit_0.register_file_0.r3_2_ ;
  wire execution_unit_0.register_file_0.r3_3_ ;
  wire execution_unit_0.register_file_0.r3_4_ ;
  wire execution_unit_0.register_file_0.r3_5_ ;
  wire execution_unit_0.register_file_0.r3_6_ ;
  wire execution_unit_0.register_file_0.r3_7_ ;
  wire execution_unit_0.register_file_0.r3_8_ ;
  wire execution_unit_0.register_file_0.r3_9_ ;
  wire execution_unit_0.register_file_0.r4_0_ ;
  wire execution_unit_0.register_file_0.r4_10_ ;
  wire execution_unit_0.register_file_0.r4_11_ ;
  wire execution_unit_0.register_file_0.r4_12_ ;
  wire execution_unit_0.register_file_0.r4_13_ ;
  wire execution_unit_0.register_file_0.r4_14_ ;
  wire execution_unit_0.register_file_0.r4_15_ ;
  wire execution_unit_0.register_file_0.r4_1_ ;
  wire execution_unit_0.register_file_0.r4_2_ ;
  wire execution_unit_0.register_file_0.r4_3_ ;
  wire execution_unit_0.register_file_0.r4_4_ ;
  wire execution_unit_0.register_file_0.r4_5_ ;
  wire execution_unit_0.register_file_0.r4_6_ ;
  wire execution_unit_0.register_file_0.r4_7_ ;
  wire execution_unit_0.register_file_0.r4_8_ ;
  wire execution_unit_0.register_file_0.r4_9_ ;
  wire execution_unit_0.register_file_0.r5_0_ ;
  wire execution_unit_0.register_file_0.r5_10_ ;
  wire execution_unit_0.register_file_0.r5_11_ ;
  wire execution_unit_0.register_file_0.r5_12_ ;
  wire execution_unit_0.register_file_0.r5_13_ ;
  wire execution_unit_0.register_file_0.r5_14_ ;
  wire execution_unit_0.register_file_0.r5_15_ ;
  wire execution_unit_0.register_file_0.r5_1_ ;
  wire execution_unit_0.register_file_0.r5_2_ ;
  wire execution_unit_0.register_file_0.r5_3_ ;
  wire execution_unit_0.register_file_0.r5_4_ ;
  wire execution_unit_0.register_file_0.r5_5_ ;
  wire execution_unit_0.register_file_0.r5_6_ ;
  wire execution_unit_0.register_file_0.r5_7_ ;
  wire execution_unit_0.register_file_0.r5_8_ ;
  wire execution_unit_0.register_file_0.r5_9_ ;
  wire execution_unit_0.register_file_0.r6_0_ ;
  wire execution_unit_0.register_file_0.r6_10_ ;
  wire execution_unit_0.register_file_0.r6_11_ ;
  wire execution_unit_0.register_file_0.r6_12_ ;
  wire execution_unit_0.register_file_0.r6_13_ ;
  wire execution_unit_0.register_file_0.r6_14_ ;
  wire execution_unit_0.register_file_0.r6_15_ ;
  wire execution_unit_0.register_file_0.r6_1_ ;
  wire execution_unit_0.register_file_0.r6_2_ ;
  wire execution_unit_0.register_file_0.r6_3_ ;
  wire execution_unit_0.register_file_0.r6_4_ ;
  wire execution_unit_0.register_file_0.r6_5_ ;
  wire execution_unit_0.register_file_0.r6_6_ ;
  wire execution_unit_0.register_file_0.r6_7_ ;
  wire execution_unit_0.register_file_0.r6_8_ ;
  wire execution_unit_0.register_file_0.r6_9_ ;
  wire execution_unit_0.register_file_0.r7_0_ ;
  wire execution_unit_0.register_file_0.r7_10_ ;
  wire execution_unit_0.register_file_0.r7_11_ ;
  wire execution_unit_0.register_file_0.r7_12_ ;
  wire execution_unit_0.register_file_0.r7_13_ ;
  wire execution_unit_0.register_file_0.r7_14_ ;
  wire execution_unit_0.register_file_0.r7_15_ ;
  wire execution_unit_0.register_file_0.r7_1_ ;
  wire execution_unit_0.register_file_0.r7_2_ ;
  wire execution_unit_0.register_file_0.r7_3_ ;
  wire execution_unit_0.register_file_0.r7_4_ ;
  wire execution_unit_0.register_file_0.r7_5_ ;
  wire execution_unit_0.register_file_0.r7_6_ ;
  wire execution_unit_0.register_file_0.r7_7_ ;
  wire execution_unit_0.register_file_0.r7_8_ ;
  wire execution_unit_0.register_file_0.r7_9_ ;
  wire execution_unit_0.register_file_0.r8_0_ ;
  wire execution_unit_0.register_file_0.r8_10_ ;
  wire execution_unit_0.register_file_0.r8_11_ ;
  wire execution_unit_0.register_file_0.r8_12_ ;
  wire execution_unit_0.register_file_0.r8_13_ ;
  wire execution_unit_0.register_file_0.r8_14_ ;
  wire execution_unit_0.register_file_0.r8_15_ ;
  wire execution_unit_0.register_file_0.r8_1_ ;
  wire execution_unit_0.register_file_0.r8_2_ ;
  wire execution_unit_0.register_file_0.r8_3_ ;
  wire execution_unit_0.register_file_0.r8_4_ ;
  wire execution_unit_0.register_file_0.r8_5_ ;
  wire execution_unit_0.register_file_0.r8_6_ ;
  wire execution_unit_0.register_file_0.r8_7_ ;
  wire execution_unit_0.register_file_0.r8_8_ ;
  wire execution_unit_0.register_file_0.r8_9_ ;
  wire execution_unit_0.register_file_0.r9_0_ ;
  wire execution_unit_0.register_file_0.r9_10_ ;
  wire execution_unit_0.register_file_0.r9_11_ ;
  wire execution_unit_0.register_file_0.r9_12_ ;
  wire execution_unit_0.register_file_0.r9_13_ ;
  wire execution_unit_0.register_file_0.r9_14_ ;
  wire execution_unit_0.register_file_0.r9_15_ ;
  wire execution_unit_0.register_file_0.r9_1_ ;
  wire execution_unit_0.register_file_0.r9_2_ ;
  wire execution_unit_0.register_file_0.r9_3_ ;
  wire execution_unit_0.register_file_0.r9_4_ ;
  wire execution_unit_0.register_file_0.r9_5_ ;
  wire execution_unit_0.register_file_0.r9_6_ ;
  wire execution_unit_0.register_file_0.r9_7_ ;
  wire execution_unit_0.register_file_0.r9_8_ ;
  wire execution_unit_0.register_file_0.r9_9_ ;
  wire fe_mb_en;
  wire fe_pmem_wait;
  wire frontend_0.e_state_nxt_0_ ;
  wire frontend_0.e_state_nxt_1_ ;
  wire frontend_0.e_state_nxt_2_ ;
  wire frontend_0.e_state_nxt_3_ ;
  wire frontend_0.exec_dext_rdy ;
  wire frontend_0.exec_dst_wr ;
  wire frontend_0.exec_jmp ;
  wire frontend_0.exec_src_wr ;
  wire frontend_0.i_state_0_ ;
  wire frontend_0.i_state_1_ ;
  wire frontend_0.i_state_2_ ;
  wire frontend_0.i_state_3_ ;
  wire frontend_0.i_state_4_ ;
  wire frontend_0.i_state_5_ ;
  wire frontend_0.inst_dest_bin_0_ ;
  wire frontend_0.inst_dest_bin_1_ ;
  wire frontend_0.inst_dest_bin_2_ ;
  wire frontend_0.inst_dest_bin_3_ ;
  wire frontend_0.inst_jmp_bin_0_ ;
  wire frontend_0.inst_jmp_bin_1_ ;
  wire frontend_0.inst_jmp_bin_2_ ;
  wire frontend_0.inst_src_bin_0_ ;
  wire frontend_0.inst_src_bin_1_ ;
  wire frontend_0.inst_src_bin_2_ ;
  wire frontend_0.inst_src_bin_3_ ;
  wire frontend_0.inst_sz_0_ ;
  wire frontend_0.inst_sz_1_ ;
  wire frontend_0.irq_addr_1_ ;
  wire frontend_0.irq_addr_2_ ;
  wire frontend_0.irq_addr_3_ ;
  wire frontend_0.irq_addr_4_ ;
  wire frontend_0.irq_addr_5_ ;
  wire frontend_0.irq_addr_6_ ;
  wire frontend_0.pmem_busy ;
  wire frontend_0.wdt_irq ;
  input irq_0_;
  input irq_10_;
  input irq_11_;
  input irq_12_;
  input irq_13_;
  input irq_1_;
  input irq_2_;
  input irq_3_;
  input irq_4_;
  input irq_5_;
  input irq_6_;
  input irq_7_;
  input irq_8_;
  input irq_9_;
  output irq_acc_0_;
  output irq_acc_10_;
  output irq_acc_11_;
  output irq_acc_12_;
  output irq_acc_13_;
  output irq_acc_1_;
  output irq_acc_2_;
  output irq_acc_3_;
  output irq_acc_4_;
  output irq_acc_5_;
  output irq_acc_6_;
  output irq_acc_7_;
  output irq_acc_8_;
  output irq_acc_9_;
  input lfxt_clk;
  output lfxt_enable;
  output lfxt_wkup;
  output mclk;
  wire mem_backbone_0.eu_mdb_in_sel_0_ ;
  wire mem_backbone_0.eu_mdb_in_sel_1_ ;
  wire mem_backbone_0.eu_per_en ;
  wire mem_backbone_0.eu_pmem_en ;
  wire mem_backbone_0.ext_mem_din_sel_0_ ;
  wire mem_backbone_0.ext_mem_din_sel_1_ ;
  wire mem_backbone_0.ext_per_en ;
  wire mem_backbone_0.ext_pmem_en ;
  wire mem_backbone_0.fe_pmem_en ;
  wire mem_backbone_0.fe_pmem_en_dly ;
  wire mem_backbone_0.per_dout_0_ ;
  wire mem_backbone_0.per_dout_10_ ;
  wire mem_backbone_0.per_dout_11_ ;
  wire mem_backbone_0.per_dout_12_ ;
  wire mem_backbone_0.per_dout_13_ ;
  wire mem_backbone_0.per_dout_14_ ;
  wire mem_backbone_0.per_dout_15_ ;
  wire mem_backbone_0.per_dout_1_ ;
  wire mem_backbone_0.per_dout_2_ ;
  wire mem_backbone_0.per_dout_3_ ;
  wire mem_backbone_0.per_dout_4_ ;
  wire mem_backbone_0.per_dout_5_ ;
  wire mem_backbone_0.per_dout_6_ ;
  wire mem_backbone_0.per_dout_7_ ;
  wire mem_backbone_0.per_dout_8_ ;
  wire mem_backbone_0.per_dout_9_ ;
  wire mem_backbone_0.per_dout_val_0_ ;
  wire mem_backbone_0.per_dout_val_10_ ;
  wire mem_backbone_0.per_dout_val_11_ ;
  wire mem_backbone_0.per_dout_val_12_ ;
  wire mem_backbone_0.per_dout_val_13_ ;
  wire mem_backbone_0.per_dout_val_14_ ;
  wire mem_backbone_0.per_dout_val_15_ ;
  wire mem_backbone_0.per_dout_val_1_ ;
  wire mem_backbone_0.per_dout_val_2_ ;
  wire mem_backbone_0.per_dout_val_3_ ;
  wire mem_backbone_0.per_dout_val_4_ ;
  wire mem_backbone_0.per_dout_val_5_ ;
  wire mem_backbone_0.per_dout_val_6_ ;
  wire mem_backbone_0.per_dout_val_7_ ;
  wire mem_backbone_0.per_dout_val_8_ ;
  wire mem_backbone_0.per_dout_val_9_ ;
  wire mem_backbone_0.pmem_dout_bckup_0_ ;
  wire mem_backbone_0.pmem_dout_bckup_1_ ;
  wire mem_backbone_0.pmem_dout_bckup_2_ ;
  wire mem_backbone_0.pmem_dout_bckup_3_ ;
  wire mem_backbone_0.pmem_dout_bckup_4_ ;
  wire mem_backbone_0.pmem_dout_bckup_5_ ;
  wire mem_backbone_0.pmem_dout_bckup_6_ ;
  wire mem_backbone_0.pmem_dout_bckup_7_ ;
  wire mem_backbone_0.pmem_dout_bckup_8_ ;
  wire mem_backbone_0.pmem_dout_bckup_sel ;
  wire multiplier_0.acc_sel ;
  wire multiplier_0.cycle_0_ ;
  wire multiplier_0.cycle_1_ ;
  wire multiplier_0.op1_0_ ;
  wire multiplier_0.op1_10_ ;
  wire multiplier_0.op1_11_ ;
  wire multiplier_0.op1_12_ ;
  wire multiplier_0.op1_13_ ;
  wire multiplier_0.op1_14_ ;
  wire multiplier_0.op1_15_ ;
  wire multiplier_0.op1_1_ ;
  wire multiplier_0.op1_2_ ;
  wire multiplier_0.op1_3_ ;
  wire multiplier_0.op1_4_ ;
  wire multiplier_0.op1_5_ ;
  wire multiplier_0.op1_6_ ;
  wire multiplier_0.op1_7_ ;
  wire multiplier_0.op1_8_ ;
  wire multiplier_0.op1_9_ ;
  wire multiplier_0.op2_0_ ;
  wire multiplier_0.op2_10_ ;
  wire multiplier_0.op2_11_ ;
  wire multiplier_0.op2_12_ ;
  wire multiplier_0.op2_13_ ;
  wire multiplier_0.op2_14_ ;
  wire multiplier_0.op2_15_ ;
  wire multiplier_0.op2_1_ ;
  wire multiplier_0.op2_2_ ;
  wire multiplier_0.op2_3_ ;
  wire multiplier_0.op2_4_ ;
  wire multiplier_0.op2_5_ ;
  wire multiplier_0.op2_6_ ;
  wire multiplier_0.op2_7_ ;
  wire multiplier_0.op2_8_ ;
  wire multiplier_0.op2_9_ ;
  wire multiplier_0.op2_wr ;
  wire multiplier_0.per_dout_0_ ;
  wire multiplier_0.per_dout_10_ ;
  wire multiplier_0.per_dout_11_ ;
  wire multiplier_0.per_dout_12_ ;
  wire multiplier_0.per_dout_13_ ;
  wire multiplier_0.per_dout_14_ ;
  wire multiplier_0.per_dout_15_ ;
  wire multiplier_0.per_dout_1_ ;
  wire multiplier_0.per_dout_2_ ;
  wire multiplier_0.per_dout_3_ ;
  wire multiplier_0.per_dout_4_ ;
  wire multiplier_0.per_dout_5_ ;
  wire multiplier_0.per_dout_6_ ;
  wire multiplier_0.per_dout_7_ ;
  wire multiplier_0.per_dout_8_ ;
  wire multiplier_0.per_dout_9_ ;
  wire multiplier_0.reshi_0_ ;
  wire multiplier_0.reshi_10_ ;
  wire multiplier_0.reshi_11_ ;
  wire multiplier_0.reshi_12_ ;
  wire multiplier_0.reshi_13_ ;
  wire multiplier_0.reshi_14_ ;
  wire multiplier_0.reshi_15_ ;
  wire multiplier_0.reshi_1_ ;
  wire multiplier_0.reshi_2_ ;
  wire multiplier_0.reshi_3_ ;
  wire multiplier_0.reshi_4_ ;
  wire multiplier_0.reshi_5_ ;
  wire multiplier_0.reshi_6_ ;
  wire multiplier_0.reshi_7_ ;
  wire multiplier_0.reshi_8_ ;
  wire multiplier_0.reshi_9_ ;
  wire multiplier_0.reslo_0_ ;
  wire multiplier_0.reslo_10_ ;
  wire multiplier_0.reslo_11_ ;
  wire multiplier_0.reslo_12_ ;
  wire multiplier_0.reslo_13_ ;
  wire multiplier_0.reslo_14_ ;
  wire multiplier_0.reslo_15_ ;
  wire multiplier_0.reslo_1_ ;
  wire multiplier_0.reslo_2_ ;
  wire multiplier_0.reslo_3_ ;
  wire multiplier_0.reslo_4_ ;
  wire multiplier_0.reslo_5_ ;
  wire multiplier_0.reslo_6_ ;
  wire multiplier_0.reslo_7_ ;
  wire multiplier_0.reslo_8_ ;
  wire multiplier_0.reslo_9_ ;
  wire multiplier_0.sign_sel ;
  wire multiplier_0.sumext_0_ ;
  wire multiplier_0.sumext_10_ ;
  input nmi;
  output per_addr_0_;
  output per_addr_10_;
  output per_addr_11_;
  output per_addr_12_;
  output per_addr_13_;
  output per_addr_1_;
  output per_addr_2_;
  output per_addr_3_;
  output per_addr_4_;
  output per_addr_5_;
  output per_addr_6_;
  output per_addr_7_;
  output per_addr_8_;
  output per_addr_9_;
  output per_din_0_;
  output per_din_10_;
  output per_din_11_;
  output per_din_12_;
  output per_din_13_;
  output per_din_14_;
  output per_din_15_;
  output per_din_1_;
  output per_din_2_;
  output per_din_3_;
  output per_din_4_;
  output per_din_5_;
  output per_din_6_;
  output per_din_7_;
  output per_din_8_;
  output per_din_9_;
  input per_dout_0_;
  input per_dout_10_;
  input per_dout_11_;
  input per_dout_12_;
  input per_dout_13_;
  input per_dout_14_;
  input per_dout_15_;
  input per_dout_1_;
  input per_dout_2_;
  input per_dout_3_;
  input per_dout_4_;
  input per_dout_5_;
  input per_dout_6_;
  input per_dout_7_;
  input per_dout_8_;
  input per_dout_9_;
  wire per_dout_sfr_0_;
  wire per_dout_sfr_10_;
  wire per_dout_sfr_11_;
  wire per_dout_sfr_12_;
  wire per_dout_sfr_13_;
  wire per_dout_sfr_14_;
  wire per_dout_sfr_15_;
  wire per_dout_sfr_1_;
  wire per_dout_sfr_2_;
  wire per_dout_sfr_3_;
  wire per_dout_sfr_4_;
  wire per_dout_sfr_5_;
  wire per_dout_sfr_6_;
  wire per_dout_sfr_7_;
  wire per_dout_sfr_8_;
  wire per_dout_sfr_9_;
  wire per_dout_wdog_0_;
  wire per_dout_wdog_11_;
  wire per_dout_wdog_1_;
  wire per_dout_wdog_2_;
  wire per_dout_wdog_3_;
  wire per_dout_wdog_4_;
  wire per_dout_wdog_5_;
  wire per_dout_wdog_6_;
  wire per_dout_wdog_7_;
  output per_en;
  output per_we_0_;
  output per_we_1_;
  output pmem_addr_0_;
  output pmem_addr_10_;
  output pmem_addr_11_;
  output pmem_addr_12_;
  output pmem_addr_13_;
  output pmem_addr_1_;
  output pmem_addr_2_;
  output pmem_addr_3_;
  output pmem_addr_4_;
  output pmem_addr_5_;
  output pmem_addr_6_;
  output pmem_addr_7_;
  output pmem_addr_8_;
  output pmem_addr_9_;
  output pmem_cen;
  output pmem_din_0_;
  output pmem_din_10_;
  output pmem_din_11_;
  output pmem_din_12_;
  output pmem_din_13_;
  output pmem_din_14_;
  output pmem_din_15_;
  output pmem_din_1_;
  output pmem_din_2_;
  output pmem_din_3_;
  output pmem_din_4_;
  output pmem_din_5_;
  output pmem_din_6_;
  output pmem_din_7_;
  output pmem_din_8_;
  output pmem_din_9_;
  input pmem_dout_0_;
  input pmem_dout_10_;
  input pmem_dout_11_;
  input pmem_dout_12_;
  input pmem_dout_13_;
  input pmem_dout_14_;
  input pmem_dout_15_;
  input pmem_dout_1_;
  input pmem_dout_2_;
  input pmem_dout_3_;
  input pmem_dout_4_;
  input pmem_dout_5_;
  input pmem_dout_6_;
  input pmem_dout_7_;
  input pmem_dout_8_;
  input pmem_dout_9_;
  output pmem_wen_0_;
  output pmem_wen_1_;
  output puc_rst;
  input reset_n;
  input scan_enable;
  input scan_mode;
  wire sfr_0.UNUSED_wdtnmies ;
  wire sfr_0.ie1_0_ ;
  wire sfr_0.ifg1_0_ ;
  wire sfr_0.wdtifg_sw_clr ;
  wire sfr_0.wdtifg_sw_set ;
  output smclk;
  output smclk_en;
  wire watchdog_0.wdtcnt_0_ ;
  wire watchdog_0.wdtcnt_10_ ;
  wire watchdog_0.wdtcnt_11_ ;
  wire watchdog_0.wdtcnt_12_ ;
  wire watchdog_0.wdtcnt_13_ ;
  wire watchdog_0.wdtcnt_14_ ;
  wire watchdog_0.wdtcnt_15_ ;
  wire watchdog_0.wdtcnt_1_ ;
  wire watchdog_0.wdtcnt_2_ ;
  wire watchdog_0.wdtcnt_3_ ;
  wire watchdog_0.wdtcnt_4_ ;
  wire watchdog_0.wdtcnt_5_ ;
  wire watchdog_0.wdtcnt_6_ ;
  wire watchdog_0.wdtcnt_7_ ;
  wire watchdog_0.wdtcnt_8_ ;
  wire watchdog_0.wdtcnt_9_ ;
  wire watchdog_0.wdtctl_0_ ;
  wire watchdog_0.wdtctl_1_ ;
  wire watchdog_0.wdtctl_2_ ;
  wire watchdog_0.wdtctl_3_ ;
  wire watchdog_0.wdtctl_4_ ;
  wire watchdog_0.wdtctl_5_ ;
  wire watchdog_0.wdtctl_7_ ;
  input wkup;
  INVX1 _06054_ (
    .A(multiplier_0.per_dout_0_ ),
    .Y(_00045_)
  );
  INVX1 _06055_ (
    .A(multiplier_0.per_dout_1_ ),
    .Y(_00046_)
  );
  INVX1 _06056_ (
    .A(multiplier_0.per_dout_2_ ),
    .Y(_00047_)
  );
  INVX1 _06057_ (
    .A(multiplier_0.per_dout_3_ ),
    .Y(_00000_)
  );
  INVX1 _06058_ (
    .A(multiplier_0.per_dout_4_ ),
    .Y(_00001_)
  );
  INVX1 _06059_ (
    .A(multiplier_0.per_dout_5_ ),
    .Y(_00002_)
  );
  INVX1 _06060_ (
    .A(multiplier_0.per_dout_6_ ),
    .Y(_00003_)
  );
  INVX1 _06061_ (
    .A(multiplier_0.per_dout_7_ ),
    .Y(_00004_)
  );
  INVX1 _06062_ (
    .A(multiplier_0.per_dout_8_ ),
    .Y(_00005_)
  );
  INVX1 _06063_ (
    .A(multiplier_0.per_dout_9_ ),
    .Y(_00006_)
  );
  INVX1 _06064_ (
    .A(multiplier_0.per_dout_10_ ),
    .Y(_00007_)
  );
  INVX1 _06065_ (
    .A(multiplier_0.per_dout_11_ ),
    .Y(_00008_)
  );
  INVX1 _06066_ (
    .A(multiplier_0.per_dout_12_ ),
    .Y(_00009_)
  );
  INVX1 _06067_ (
    .A(multiplier_0.per_dout_13_ ),
    .Y(_00010_)
  );
  INVX1 _06068_ (
    .A(multiplier_0.per_dout_14_ ),
    .Y(_00011_)
  );
  INVX1 _06069_ (
    .A(multiplier_0.per_dout_15_ ),
    .Y(_00012_)
  );
  NOR2X1 _06070_ (
    .A(clock_module_0.bcsctl2_rd_0_ ),
    .B(per_dout_0_),
    .Y(_00013_)
  );
  NOR2X1 _06071_ (
    .A(per_dout_sfr_0_),
    .B(per_dout_wdog_0_),
    .Y(_00014_)
  );
  NAND3X1 _06072_ (
    .A(_00045_),
    .B(_00013_),
    .C(_00014_),
    .Y(mem_backbone_0.per_dout_0_ )
  );
  NOR2X1 _06073_ (
    .A(clock_module_0.bcsctl2_rd_1_ ),
    .B(per_dout_1_),
    .Y(_00015_)
  );
  NOR2X1 _06074_ (
    .A(per_dout_sfr_1_),
    .B(per_dout_wdog_1_),
    .Y(_00016_)
  );
  NAND3X1 _06075_ (
    .A(_00046_),
    .B(_00015_),
    .C(_00016_),
    .Y(mem_backbone_0.per_dout_1_ )
  );
  NOR2X1 _06076_ (
    .A(clock_module_0.bcsctl2_rd_2_ ),
    .B(per_dout_2_),
    .Y(_00017_)
  );
  NOR2X1 _06077_ (
    .A(per_dout_sfr_2_),
    .B(per_dout_wdog_2_),
    .Y(_00018_)
  );
  NAND3X1 _06078_ (
    .A(_00047_),
    .B(_00017_),
    .C(_00018_),
    .Y(mem_backbone_0.per_dout_2_ )
  );
  NOR2X1 _06079_ (
    .A(clock_module_0.bcsctl2_rd_3_ ),
    .B(per_dout_3_),
    .Y(_00019_)
  );
  NOR2X1 _06080_ (
    .A(per_dout_sfr_3_),
    .B(per_dout_wdog_3_),
    .Y(_00020_)
  );
  NAND3X1 _06081_ (
    .A(_00000_),
    .B(_00019_),
    .C(_00020_),
    .Y(mem_backbone_0.per_dout_3_ )
  );
  NOR2X1 _06082_ (
    .A(clock_module_0.bcsctl2_rd_4_ ),
    .B(per_dout_4_),
    .Y(_00021_)
  );
  NOR2X1 _06083_ (
    .A(per_dout_sfr_4_),
    .B(per_dout_wdog_4_),
    .Y(_00022_)
  );
  NAND3X1 _06084_ (
    .A(_00001_),
    .B(_00021_),
    .C(_00022_),
    .Y(mem_backbone_0.per_dout_4_ )
  );
  NOR2X1 _06085_ (
    .A(clock_module_0.bcsctl2_rd_5_ ),
    .B(per_dout_5_),
    .Y(_00023_)
  );
  NOR2X1 _06086_ (
    .A(per_dout_sfr_5_),
    .B(per_dout_wdog_5_),
    .Y(_00024_)
  );
  NAND3X1 _06087_ (
    .A(_00002_),
    .B(_00023_),
    .C(_00024_),
    .Y(mem_backbone_0.per_dout_5_ )
  );
  NOR2X1 _06088_ (
    .A(clock_module_0.bcsctl2_rd_6_ ),
    .B(per_dout_6_),
    .Y(_00025_)
  );
  NOR2X1 _06089_ (
    .A(per_dout_sfr_6_),
    .B(per_dout_wdog_6_),
    .Y(_00026_)
  );
  NAND3X1 _06090_ (
    .A(_00003_),
    .B(_00025_),
    .C(_00026_),
    .Y(mem_backbone_0.per_dout_6_ )
  );
  NOR2X1 _06091_ (
    .A(clock_module_0.bcsctl2_rd_7_ ),
    .B(per_dout_7_),
    .Y(_00027_)
  );
  NOR2X1 _06092_ (
    .A(per_dout_sfr_7_),
    .B(per_dout_wdog_7_),
    .Y(_00028_)
  );
  NAND3X1 _06093_ (
    .A(_00004_),
    .B(_00027_),
    .C(_00028_),
    .Y(mem_backbone_0.per_dout_7_ )
  );
  NOR2X1 _06094_ (
    .A(clock_module_0.bcsctl1_rd_8_ ),
    .B(per_dout_8_),
    .Y(_00029_)
  );
  NOR2X1 _06095_ (
    .A(per_dout_sfr_8_),
    .B(per_dout_wdog_11_),
    .Y(_00030_)
  );
  NAND3X1 _06096_ (
    .A(_00005_),
    .B(_00029_),
    .C(_00030_),
    .Y(mem_backbone_0.per_dout_8_ )
  );
  NOR2X1 _06097_ (
    .A(clock_module_0.bcsctl1_rd_9_ ),
    .B(per_dout_9_),
    .Y(_00031_)
  );
  NOR2X1 _06098_ (
    .A(per_dout_sfr_9_),
    .B(1'h0),
    .Y(_00032_)
  );
  NAND3X1 _06099_ (
    .A(_00006_),
    .B(_00031_),
    .C(_00032_),
    .Y(mem_backbone_0.per_dout_9_ )
  );
  NOR2X1 _06100_ (
    .A(clock_module_0.bcsctl1_rd_10_ ),
    .B(per_dout_10_),
    .Y(_00033_)
  );
  NOR2X1 _06101_ (
    .A(per_dout_sfr_10_),
    .B(1'h0),
    .Y(_00034_)
  );
  NAND3X1 _06102_ (
    .A(_00007_),
    .B(_00033_),
    .C(_00034_),
    .Y(mem_backbone_0.per_dout_10_ )
  );
  NOR2X1 _06103_ (
    .A(clock_module_0.bcsctl1_rd_11_ ),
    .B(per_dout_11_),
    .Y(_00035_)
  );
  NOR2X1 _06104_ (
    .A(per_dout_sfr_11_),
    .B(per_dout_wdog_11_),
    .Y(_00036_)
  );
  NAND3X1 _06105_ (
    .A(_00008_),
    .B(_00035_),
    .C(_00036_),
    .Y(mem_backbone_0.per_dout_11_ )
  );
  NOR2X1 _06106_ (
    .A(clock_module_0.bcsctl1_rd_12_ ),
    .B(per_dout_12_),
    .Y(_00037_)
  );
  NOR2X1 _06107_ (
    .A(per_dout_sfr_12_),
    .B(1'h0),
    .Y(_00038_)
  );
  NAND3X1 _06108_ (
    .A(_00009_),
    .B(_00037_),
    .C(_00038_),
    .Y(mem_backbone_0.per_dout_12_ )
  );
  NOR2X1 _06109_ (
    .A(clock_module_0.bcsctl1_rd_13_ ),
    .B(per_dout_13_),
    .Y(_00039_)
  );
  NOR2X1 _06110_ (
    .A(per_dout_sfr_13_),
    .B(per_dout_wdog_11_),
    .Y(_00040_)
  );
  NAND3X1 _06111_ (
    .A(_00010_),
    .B(_00039_),
    .C(_00040_),
    .Y(mem_backbone_0.per_dout_13_ )
  );
  NOR2X1 _06112_ (
    .A(clock_module_0.bcsctl1_rd_14_ ),
    .B(per_dout_14_),
    .Y(_00041_)
  );
  NOR2X1 _06113_ (
    .A(per_dout_sfr_14_),
    .B(per_dout_wdog_11_),
    .Y(_00042_)
  );
  NAND3X1 _06114_ (
    .A(_00011_),
    .B(_00041_),
    .C(_00042_),
    .Y(mem_backbone_0.per_dout_14_ )
  );
  NOR2X1 _06115_ (
    .A(clock_module_0.bcsctl1_rd_15_ ),
    .B(per_dout_15_),
    .Y(_00043_)
  );
  NOR2X1 _06116_ (
    .A(per_dout_sfr_15_),
    .B(1'h0),
    .Y(_00044_)
  );
  NAND3X1 _06117_ (
    .A(_00012_),
    .B(_00043_),
    .C(_00044_),
    .Y(mem_backbone_0.per_dout_15_ )
  );
  BUFX2 _06118_ (
    .A(dco_clk),
    .Y(aclk)
  );
  BUFX2 _06119_ (
    .A(_00048_),
    .Y(aclk_en)
  );
  BUFX2 _06120_ (
    .A(_00049_),
    .Y(dbg_freeze)
  );
  BUFX2 _06121_ (
    .A(_00050_),
    .Y(dbg_i2c_sda_out)
  );
  BUFX2 _06122_ (
    .A(1'h1),
    .Y(dbg_uart_txd)
  );
  BUFX2 _06123_ (
    .A(1'h1),
    .Y(dco_enable)
  );
  BUFX2 _06124_ (
    .A(1'h1),
    .Y(dco_wkup)
  );
  BUFX2 _06125_ (
    .A(1'h0),
    .Y(dma_dout_0_)
  );
  BUFX2 _06126_ (
    .A(1'h0),
    .Y(dma_dout_10_)
  );
  BUFX2 _06127_ (
    .A(1'h0),
    .Y(dma_dout_11_)
  );
  BUFX2 _06128_ (
    .A(1'h0),
    .Y(dma_dout_12_)
  );
  BUFX2 _06129_ (
    .A(1'h0),
    .Y(dma_dout_13_)
  );
  BUFX2 _06130_ (
    .A(1'h0),
    .Y(dma_dout_14_)
  );
  BUFX2 _06131_ (
    .A(1'h0),
    .Y(dma_dout_15_)
  );
  BUFX2 _06132_ (
    .A(1'h0),
    .Y(dma_dout_1_)
  );
  BUFX2 _06133_ (
    .A(1'h0),
    .Y(dma_dout_2_)
  );
  BUFX2 _06134_ (
    .A(1'h0),
    .Y(dma_dout_3_)
  );
  BUFX2 _06135_ (
    .A(1'h0),
    .Y(dma_dout_4_)
  );
  BUFX2 _06136_ (
    .A(1'h0),
    .Y(dma_dout_5_)
  );
  BUFX2 _06137_ (
    .A(1'h0),
    .Y(dma_dout_6_)
  );
  BUFX2 _06138_ (
    .A(1'h0),
    .Y(dma_dout_7_)
  );
  BUFX2 _06139_ (
    .A(1'h0),
    .Y(dma_dout_8_)
  );
  BUFX2 _06140_ (
    .A(1'h0),
    .Y(dma_dout_9_)
  );
  BUFX2 _06141_ (
    .A(1'h1),
    .Y(dma_ready)
  );
  BUFX2 _06142_ (
    .A(1'h1),
    .Y(dma_resp)
  );
  BUFX2 _06143_ (
    .A(_00051_),
    .Y(dmem_addr_0_)
  );
  BUFX2 _06144_ (
    .A(_00052_),
    .Y(dmem_addr_10_)
  );
  BUFX2 _06145_ (
    .A(_00053_),
    .Y(dmem_addr_11_)
  );
  BUFX2 _06146_ (
    .A(_00054_),
    .Y(dmem_addr_12_)
  );
  BUFX2 _06147_ (
    .A(_00055_),
    .Y(dmem_addr_1_)
  );
  BUFX2 _06148_ (
    .A(_00056_),
    .Y(dmem_addr_2_)
  );
  BUFX2 _06149_ (
    .A(_00057_),
    .Y(dmem_addr_3_)
  );
  BUFX2 _06150_ (
    .A(_00058_),
    .Y(dmem_addr_4_)
  );
  BUFX2 _06151_ (
    .A(_00059_),
    .Y(dmem_addr_5_)
  );
  BUFX2 _06152_ (
    .A(_00060_),
    .Y(dmem_addr_6_)
  );
  BUFX2 _06153_ (
    .A(_00061_),
    .Y(dmem_addr_7_)
  );
  BUFX2 _06154_ (
    .A(_00062_),
    .Y(dmem_addr_8_)
  );
  BUFX2 _06155_ (
    .A(_00063_),
    .Y(dmem_addr_9_)
  );
  BUFX2 _06156_ (
    .A(_00064_),
    .Y(dmem_cen)
  );
  BUFX2 _06157_ (
    .A(_00065_),
    .Y(dmem_din_0_)
  );
  BUFX2 _06158_ (
    .A(_00066_),
    .Y(dmem_din_10_)
  );
  BUFX2 _06159_ (
    .A(_00067_),
    .Y(dmem_din_11_)
  );
  BUFX2 _06160_ (
    .A(_00068_),
    .Y(dmem_din_12_)
  );
  BUFX2 _06161_ (
    .A(_00069_),
    .Y(dmem_din_13_)
  );
  BUFX2 _06162_ (
    .A(_00070_),
    .Y(dmem_din_14_)
  );
  BUFX2 _06163_ (
    .A(_00071_),
    .Y(dmem_din_15_)
  );
  BUFX2 _06164_ (
    .A(_00072_),
    .Y(dmem_din_1_)
  );
  BUFX2 _06165_ (
    .A(_00073_),
    .Y(dmem_din_2_)
  );
  BUFX2 _06166_ (
    .A(_00074_),
    .Y(dmem_din_3_)
  );
  BUFX2 _06167_ (
    .A(_00075_),
    .Y(dmem_din_4_)
  );
  BUFX2 _06168_ (
    .A(_00076_),
    .Y(dmem_din_5_)
  );
  BUFX2 _06169_ (
    .A(_00077_),
    .Y(dmem_din_6_)
  );
  BUFX2 _06170_ (
    .A(_00078_),
    .Y(dmem_din_7_)
  );
  BUFX2 _06171_ (
    .A(_00079_),
    .Y(dmem_din_8_)
  );
  BUFX2 _06172_ (
    .A(_00080_),
    .Y(dmem_din_9_)
  );
  BUFX2 _06173_ (
    .A(_00081_),
    .Y(dmem_wen_0_)
  );
  BUFX2 _06174_ (
    .A(_00082_),
    .Y(dmem_wen_1_)
  );
  BUFX2 _06175_ (
    .A(_00083_),
    .Y(irq_acc_0_)
  );
  BUFX2 _06176_ (
    .A(_00084_),
    .Y(irq_acc_10_)
  );
  BUFX2 _06177_ (
    .A(_00085_),
    .Y(irq_acc_11_)
  );
  BUFX2 _06178_ (
    .A(_00086_),
    .Y(irq_acc_12_)
  );
  BUFX2 _06179_ (
    .A(_00087_),
    .Y(irq_acc_13_)
  );
  BUFX2 _06180_ (
    .A(_00088_),
    .Y(irq_acc_1_)
  );
  BUFX2 _06181_ (
    .A(_00089_),
    .Y(irq_acc_2_)
  );
  BUFX2 _06182_ (
    .A(_00090_),
    .Y(irq_acc_3_)
  );
  BUFX2 _06183_ (
    .A(_00091_),
    .Y(irq_acc_4_)
  );
  BUFX2 _06184_ (
    .A(_00092_),
    .Y(irq_acc_5_)
  );
  BUFX2 _06185_ (
    .A(_00093_),
    .Y(irq_acc_6_)
  );
  BUFX2 _06186_ (
    .A(_00094_),
    .Y(irq_acc_7_)
  );
  BUFX2 _06187_ (
    .A(_00095_),
    .Y(irq_acc_8_)
  );
  BUFX2 _06188_ (
    .A(_00096_),
    .Y(irq_acc_9_)
  );
  BUFX2 _06189_ (
    .A(1'h1),
    .Y(lfxt_enable)
  );
  BUFX2 _06190_ (
    .A(1'h0),
    .Y(lfxt_wkup)
  );
  BUFX2 _06191_ (
    .A(dco_clk),
    .Y(mclk)
  );
  BUFX2 _06192_ (
    .A(_00097_),
    .Y(per_addr_0_)
  );
  BUFX2 _06193_ (
    .A(_00098_),
    .Y(per_addr_10_)
  );
  BUFX2 _06194_ (
    .A(_00099_),
    .Y(per_addr_11_)
  );
  BUFX2 _06195_ (
    .A(_00100_),
    .Y(per_addr_12_)
  );
  BUFX2 _06196_ (
    .A(1'h0),
    .Y(per_addr_13_)
  );
  BUFX2 _06197_ (
    .A(_00101_),
    .Y(per_addr_1_)
  );
  BUFX2 _06198_ (
    .A(_00102_),
    .Y(per_addr_2_)
  );
  BUFX2 _06199_ (
    .A(_00103_),
    .Y(per_addr_3_)
  );
  BUFX2 _06200_ (
    .A(_00104_),
    .Y(per_addr_4_)
  );
  BUFX2 _06201_ (
    .A(_00105_),
    .Y(per_addr_5_)
  );
  BUFX2 _06202_ (
    .A(_00106_),
    .Y(per_addr_6_)
  );
  BUFX2 _06203_ (
    .A(_00107_),
    .Y(per_addr_7_)
  );
  BUFX2 _06204_ (
    .A(_00108_),
    .Y(per_addr_8_)
  );
  BUFX2 _06205_ (
    .A(_00109_),
    .Y(per_addr_9_)
  );
  BUFX2 _06206_ (
    .A(_00110_),
    .Y(per_din_0_)
  );
  BUFX2 _06207_ (
    .A(_00111_),
    .Y(per_din_10_)
  );
  BUFX2 _06208_ (
    .A(_00112_),
    .Y(per_din_11_)
  );
  BUFX2 _06209_ (
    .A(_00113_),
    .Y(per_din_12_)
  );
  BUFX2 _06210_ (
    .A(_00114_),
    .Y(per_din_13_)
  );
  BUFX2 _06211_ (
    .A(_00115_),
    .Y(per_din_14_)
  );
  BUFX2 _06212_ (
    .A(_00116_),
    .Y(per_din_15_)
  );
  BUFX2 _06213_ (
    .A(_00117_),
    .Y(per_din_1_)
  );
  BUFX2 _06214_ (
    .A(_00118_),
    .Y(per_din_2_)
  );
  BUFX2 _06215_ (
    .A(_00119_),
    .Y(per_din_3_)
  );
  BUFX2 _06216_ (
    .A(_00120_),
    .Y(per_din_4_)
  );
  BUFX2 _06217_ (
    .A(_00121_),
    .Y(per_din_5_)
  );
  BUFX2 _06218_ (
    .A(_00122_),
    .Y(per_din_6_)
  );
  BUFX2 _06219_ (
    .A(_00123_),
    .Y(per_din_7_)
  );
  BUFX2 _06220_ (
    .A(_00124_),
    .Y(per_din_8_)
  );
  BUFX2 _06221_ (
    .A(_00125_),
    .Y(per_din_9_)
  );
  BUFX2 _06222_ (
    .A(_00126_),
    .Y(per_en)
  );
  BUFX2 _06223_ (
    .A(_00127_),
    .Y(per_we_0_)
  );
  BUFX2 _06224_ (
    .A(_00128_),
    .Y(per_we_1_)
  );
  BUFX2 _06225_ (
    .A(_00129_),
    .Y(pmem_addr_0_)
  );
  BUFX2 _06226_ (
    .A(_00130_),
    .Y(pmem_addr_10_)
  );
  BUFX2 _06227_ (
    .A(_00131_),
    .Y(pmem_addr_11_)
  );
  BUFX2 _06228_ (
    .A(_00132_),
    .Y(pmem_addr_12_)
  );
  BUFX2 _06229_ (
    .A(_00133_),
    .Y(pmem_addr_13_)
  );
  BUFX2 _06230_ (
    .A(_00134_),
    .Y(pmem_addr_1_)
  );
  BUFX2 _06231_ (
    .A(_00135_),
    .Y(pmem_addr_2_)
  );
  BUFX2 _06232_ (
    .A(_00136_),
    .Y(pmem_addr_3_)
  );
  BUFX2 _06233_ (
    .A(_00137_),
    .Y(pmem_addr_4_)
  );
  BUFX2 _06234_ (
    .A(_00138_),
    .Y(pmem_addr_5_)
  );
  BUFX2 _06235_ (
    .A(_00139_),
    .Y(pmem_addr_6_)
  );
  BUFX2 _06236_ (
    .A(_00140_),
    .Y(pmem_addr_7_)
  );
  BUFX2 _06237_ (
    .A(_00141_),
    .Y(pmem_addr_8_)
  );
  BUFX2 _06238_ (
    .A(_00142_),
    .Y(pmem_addr_9_)
  );
  BUFX2 _06239_ (
    .A(_00143_),
    .Y(pmem_cen)
  );
  BUFX2 _06240_ (
    .A(_00144_),
    .Y(pmem_din_0_)
  );
  BUFX2 _06241_ (
    .A(_00145_),
    .Y(pmem_din_10_)
  );
  BUFX2 _06242_ (
    .A(_00146_),
    .Y(pmem_din_11_)
  );
  BUFX2 _06243_ (
    .A(_00147_),
    .Y(pmem_din_12_)
  );
  BUFX2 _06244_ (
    .A(_00148_),
    .Y(pmem_din_13_)
  );
  BUFX2 _06245_ (
    .A(_00149_),
    .Y(pmem_din_14_)
  );
  BUFX2 _06246_ (
    .A(_00150_),
    .Y(pmem_din_15_)
  );
  BUFX2 _06247_ (
    .A(_00151_),
    .Y(pmem_din_1_)
  );
  BUFX2 _06248_ (
    .A(_00152_),
    .Y(pmem_din_2_)
  );
  BUFX2 _06249_ (
    .A(_00153_),
    .Y(pmem_din_3_)
  );
  BUFX2 _06250_ (
    .A(_00154_),
    .Y(pmem_din_4_)
  );
  BUFX2 _06251_ (
    .A(_00155_),
    .Y(pmem_din_5_)
  );
  BUFX2 _06252_ (
    .A(_00156_),
    .Y(pmem_din_6_)
  );
  BUFX2 _06253_ (
    .A(_00157_),
    .Y(pmem_din_7_)
  );
  BUFX2 _06254_ (
    .A(_00158_),
    .Y(pmem_din_8_)
  );
  BUFX2 _06255_ (
    .A(_00159_),
    .Y(pmem_din_9_)
  );
  BUFX2 _06256_ (
    .A(_00160_),
    .Y(pmem_wen_0_)
  );
  BUFX2 _06257_ (
    .A(_00161_),
    .Y(pmem_wen_1_)
  );
  BUFX2 _06258_ (
    .A(_00162_),
    .Y(puc_rst)
  );
  BUFX2 _06259_ (
    .A(dco_clk),
    .Y(smclk)
  );
  BUFX2 _06260_ (
    .A(_00163_),
    .Y(smclk_en)
  );
  INVX1 _06261_ (
    .A(reset_n),
    .Y(clock_module_0.por_a )
  );
  INVX1 _06262_ (
    .A(_00104_),
    .Y(_00189_)
  );
  INVX1 _06263_ (
    .A(_00106_),
    .Y(_00190_)
  );
  INVX1 _06264_ (
    .A(_00100_),
    .Y(_00191_)
  );
  INVX1 _06265_ (
    .A(clock_module_0.bcsctl1_4_ ),
    .Y(_00192_)
  );
  INVX1 _06266_ (
    .A(clock_module_0.lfxt_clk_s ),
    .Y(_00193_)
  );
  INVX1 _06267_ (
    .A(clock_module_0.bcsctl2_1_ ),
    .Y(_00194_)
  );
  INVX1 _06268_ (
    .A(clock_module_0.bcsctl2_3_ ),
    .Y(_00195_)
  );
  INVX1 _06269_ (
    .A(clock_module_0.scg1 ),
    .Y(_00196_)
  );
  INVX1 _06270_ (
    .A(dbg_en),
    .Y(clock_module_0.dbg_rst_nxt )
  );
  INVX1 _06271_ (
    .A(clock_module_0.puc_noscan_n ),
    .Y(_00162_)
  );
  INVX1 _06272_ (
    .A(clock_module_0.por ),
    .Y(_00188_)
  );
  NOR2X1 _06273_ (
    .A(_00099_),
    .B(1'h0),
    .Y(_00197_)
  );
  NAND3X1 _06274_ (
    .A(_00191_),
    .B(_00126_),
    .C(_00197_),
    .Y(_00198_)
  );
  INVX1 _06275_ (
    .A(_00198_),
    .Y(_00199_)
  );
  NOR2X1 _06276_ (
    .A(_00108_),
    .B(_00107_),
    .Y(_00200_)
  );
  NOR2X1 _06277_ (
    .A(_00098_),
    .B(_00109_),
    .Y(_00201_)
  );
  NAND2X1 _06278_ (
    .A(_00200_),
    .B(_00201_),
    .Y(_00202_)
  );
  NAND2X1 _06279_ (
    .A(_00189_),
    .B(_00103_),
    .Y(_00203_)
  );
  NAND2X1 _06280_ (
    .A(_00190_),
    .B(_00105_),
    .Y(_00204_)
  );
  NOR3X1 _06281_ (
    .A(_00202_),
    .B(_00203_),
    .C(_00204_),
    .Y(_00205_)
  );
  NAND2X1 _06282_ (
    .A(_00101_),
    .B(_00097_),
    .Y(_00206_)
  );
  NOR2X1 _06283_ (
    .A(_00102_),
    .B(_00206_),
    .Y(_00207_)
  );
  NOR2X1 _06284_ (
    .A(_00108_),
    .B(_00109_),
    .Y(_00208_)
  );
  NAND3X1 _06285_ (
    .A(_00189_),
    .B(_00190_),
    .C(_00208_),
    .Y(_00209_)
  );
  NOR2X1 _06286_ (
    .A(_00107_),
    .B(_00098_),
    .Y(_00210_)
  );
  NAND3X1 _06287_ (
    .A(_00103_),
    .B(_00105_),
    .C(_00210_),
    .Y(_00211_)
  );
  NOR3X1 _06288_ (
    .A(_00198_),
    .B(_00209_),
    .C(_00211_),
    .Y(_00212_)
  );
  NAND3X1 _06289_ (
    .A(_00128_),
    .B(_00207_),
    .C(_00212_),
    .Y(_00213_)
  );
  AND2X1 _06290_ (
    .A(clock_module_0.bcsctl1_0_ ),
    .B(_00213_),
    .Y(_00168_)
  );
  AND2X1 _06291_ (
    .A(clock_module_0.bcsctl1_1_ ),
    .B(_00213_),
    .Y(_00169_)
  );
  AND2X1 _06292_ (
    .A(clock_module_0.bcsctl1_2_ ),
    .B(_00213_),
    .Y(_00170_)
  );
  AND2X1 _06293_ (
    .A(clock_module_0.bcsctl1_3_ ),
    .B(_00213_),
    .Y(_00171_)
  );
  MUX2X1 _06294_ (
    .A(clock_module_0.bcsctl1_4_ ),
    .B(_00113_),
    .S(_00213_),
    .Y(_00214_)
  );
  INVX1 _06295_ (
    .A(_00214_),
    .Y(_00172_)
  );
  MUX2X1 _06296_ (
    .A(clock_module_0.bcsctl1_5_ ),
    .B(_00114_),
    .S(_00213_),
    .Y(_00215_)
  );
  INVX1 _06297_ (
    .A(_00215_),
    .Y(_00173_)
  );
  AND2X1 _06298_ (
    .A(clock_module_0.bcsctl1_6_ ),
    .B(_00213_),
    .Y(_00174_)
  );
  AND2X1 _06299_ (
    .A(clock_module_0.bcsctl1_7_ ),
    .B(_00213_),
    .Y(_00175_)
  );
  NOR2X1 _06300_ (
    .A(clock_module_0.bcsctl1_4_ ),
    .B(clock_module_0.bcsctl1_5_ ),
    .Y(_00216_)
  );
  NAND2X1 _06301_ (
    .A(clock_module_0.bcsctl1_1_ ),
    .B(1'h1),
    .Y(_00217_)
  );
  NAND2X1 _06302_ (
    .A(clock_module_0.oscoff ),
    .B(_00217_),
    .Y(_00218_)
  );
  NOR2X1 _06303_ (
    .A(clock_module_0.lfxt_clk_dly ),
    .B(_00193_),
    .Y(_00219_)
  );
  NAND2X1 _06304_ (
    .A(_00218_),
    .B(_00219_),
    .Y(_00220_)
  );
  NOR2X1 _06305_ (
    .A(_00216_),
    .B(_00220_),
    .Y(_00221_)
  );
  NAND2X1 _06306_ (
    .A(clock_module_0.aclk_div_0_ ),
    .B(_00221_),
    .Y(_00222_)
  );
  XOR2X1 _06307_ (
    .A(clock_module_0.aclk_div_0_ ),
    .B(_00221_),
    .Y(_00164_)
  );
  NAND3X1 _06308_ (
    .A(clock_module_0.aclk_div_0_ ),
    .B(clock_module_0.aclk_div_1_ ),
    .C(_00221_),
    .Y(_00223_)
  );
  XNOR2X1 _06309_ (
    .A(clock_module_0.aclk_div_1_ ),
    .B(_00222_),
    .Y(_00165_)
  );
  XNOR2X1 _06310_ (
    .A(clock_module_0.aclk_div_2_ ),
    .B(_00223_),
    .Y(_00166_)
  );
  AOI21X1 _06311_ (
    .A(clock_module_0.bcsctl1_3_ ),
    .B(1'h1),
    .C(_00196_),
    .Y(_00224_)
  );
  AOI21X1 _06312_ (
    .A(_00218_),
    .B(_00219_),
    .C(_00195_),
    .Y(_00225_)
  );
  NOR2X1 _06313_ (
    .A(_00224_),
    .B(_00225_),
    .Y(_00226_)
  );
  NOR2X1 _06314_ (
    .A(clock_module_0.bcsctl2_1_ ),
    .B(clock_module_0.bcsctl2_2_ ),
    .Y(_00227_)
  );
  NOR3X1 _06315_ (
    .A(_00224_),
    .B(_00225_),
    .C(_00227_),
    .Y(_00228_)
  );
  AND2X1 _06316_ (
    .A(clock_module_0.smclk_div_0_ ),
    .B(_00228_),
    .Y(_00229_)
  );
  NOR2X1 _06317_ (
    .A(clock_module_0.smclk_div_0_ ),
    .B(_00228_),
    .Y(_00230_)
  );
  NOR2X1 _06318_ (
    .A(_00229_),
    .B(_00230_),
    .Y(_00184_)
  );
  NAND3X1 _06319_ (
    .A(clock_module_0.smclk_div_0_ ),
    .B(clock_module_0.smclk_div_1_ ),
    .C(_00228_),
    .Y(_00231_)
  );
  XOR2X1 _06320_ (
    .A(clock_module_0.smclk_div_1_ ),
    .B(_00229_),
    .Y(_00185_)
  );
  XNOR2X1 _06321_ (
    .A(clock_module_0.smclk_div_2_ ),
    .B(_00231_),
    .Y(_00186_)
  );
  NOR2X1 _06322_ (
    .A(_00101_),
    .B(_00097_),
    .Y(_00232_)
  );
  AND2X1 _06323_ (
    .A(_00102_),
    .B(_00232_),
    .Y(_00233_)
  );
  NAND2X1 _06324_ (
    .A(_00102_),
    .B(_00232_),
    .Y(_00234_)
  );
  NAND3X1 _06325_ (
    .A(_00127_),
    .B(_00212_),
    .C(_00233_),
    .Y(_00235_)
  );
  AND2X1 _06326_ (
    .A(clock_module_0.bcsctl2_0_ ),
    .B(_00235_),
    .Y(_00176_)
  );
  MUX2X1 _06327_ (
    .A(clock_module_0.bcsctl2_1_ ),
    .B(_00117_),
    .S(_00235_),
    .Y(_00236_)
  );
  INVX1 _06328_ (
    .A(_00236_),
    .Y(_00177_)
  );
  MUX2X1 _06329_ (
    .A(clock_module_0.bcsctl2_2_ ),
    .B(_00118_),
    .S(_00235_),
    .Y(_00237_)
  );
  INVX1 _06330_ (
    .A(_00237_),
    .Y(_00178_)
  );
  MUX2X1 _06331_ (
    .A(clock_module_0.bcsctl2_3_ ),
    .B(_00119_),
    .S(_00235_),
    .Y(_00238_)
  );
  INVX1 _06332_ (
    .A(_00238_),
    .Y(_00179_)
  );
  AND2X1 _06333_ (
    .A(clock_module_0.bcsctl2_4_ ),
    .B(_00235_),
    .Y(_00180_)
  );
  AND2X1 _06334_ (
    .A(clock_module_0.bcsctl2_5_ ),
    .B(_00235_),
    .Y(_00181_)
  );
  AND2X1 _06335_ (
    .A(clock_module_0.bcsctl2_6_ ),
    .B(_00235_),
    .Y(_00182_)
  );
  AND2X1 _06336_ (
    .A(clock_module_0.bcsctl2_7_ ),
    .B(_00235_),
    .Y(_00183_)
  );
  NOR2X1 _06337_ (
    .A(clock_module_0.dbg_rst_nxt ),
    .B(clock_module_0.puc_noscan_n ),
    .Y(_00239_)
  );
  AOI21X1 _06338_ (
    .A(clock_module_0.dbg_rst ),
    .B(_00239_),
    .C(clock_module_0.dbg_cpu_reset ),
    .Y(clock_module_0.sync_cell_puc.data_in )
  );
  NOR2X1 _06339_ (
    .A(_00128_),
    .B(_00127_),
    .Y(_00240_)
  );
  NAND3X1 _06340_ (
    .A(_00199_),
    .B(_00205_),
    .C(_00240_),
    .Y(_00241_)
  );
  NOR3X1 _06341_ (
    .A(_00102_),
    .B(_00206_),
    .C(_00241_),
    .Y(_00242_)
  );
  AND2X1 _06342_ (
    .A(clock_module_0.bcsctl1_0_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_8_ )
  );
  AND2X1 _06343_ (
    .A(clock_module_0.bcsctl1_1_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_9_ )
  );
  AND2X1 _06344_ (
    .A(clock_module_0.bcsctl1_2_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_10_ )
  );
  AND2X1 _06345_ (
    .A(clock_module_0.bcsctl1_3_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_11_ )
  );
  AND2X1 _06346_ (
    .A(clock_module_0.bcsctl1_4_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_12_ )
  );
  AND2X1 _06347_ (
    .A(clock_module_0.bcsctl1_5_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_13_ )
  );
  AND2X1 _06348_ (
    .A(clock_module_0.bcsctl1_6_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_14_ )
  );
  AND2X1 _06349_ (
    .A(clock_module_0.bcsctl1_7_ ),
    .B(_00242_),
    .Y(clock_module_0.bcsctl1_rd_15_ )
  );
  NOR2X1 _06350_ (
    .A(_00234_),
    .B(_00241_),
    .Y(_00243_)
  );
  AND2X1 _06351_ (
    .A(clock_module_0.bcsctl2_0_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_0_ )
  );
  AND2X1 _06352_ (
    .A(clock_module_0.bcsctl2_1_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_1_ )
  );
  AND2X1 _06353_ (
    .A(clock_module_0.bcsctl2_2_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_2_ )
  );
  AND2X1 _06354_ (
    .A(clock_module_0.bcsctl2_3_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_3_ )
  );
  AND2X1 _06355_ (
    .A(clock_module_0.bcsctl2_4_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_4_ )
  );
  AND2X1 _06356_ (
    .A(clock_module_0.bcsctl2_5_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_5_ )
  );
  AND2X1 _06357_ (
    .A(clock_module_0.bcsctl2_6_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_6_ )
  );
  AND2X1 _06358_ (
    .A(clock_module_0.bcsctl2_7_ ),
    .B(_00243_),
    .Y(clock_module_0.bcsctl2_rd_7_ )
  );
  OAI21X1 _06359_ (
    .A(_00192_),
    .B(clock_module_0.aclk_div_2_ ),
    .C(clock_module_0.aclk_div_1_ ),
    .Y(_00244_)
  );
  OAI21X1 _06360_ (
    .A(clock_module_0.aclk_div_0_ ),
    .B(_00216_),
    .C(cpu_en),
    .Y(_00245_)
  );
  OR2X1 _06361_ (
    .A(_00220_),
    .B(_00245_),
    .Y(_00246_)
  );
  AOI21X1 _06362_ (
    .A(clock_module_0.bcsctl1_5_ ),
    .B(_00244_),
    .C(_00246_),
    .Y(_00167_)
  );
  OAI21X1 _06363_ (
    .A(_00194_),
    .B(clock_module_0.smclk_div_2_ ),
    .C(clock_module_0.smclk_div_1_ ),
    .Y(_00247_)
  );
  OAI21X1 _06364_ (
    .A(clock_module_0.smclk_div_0_ ),
    .B(_00227_),
    .C(cpu_en),
    .Y(_00248_)
  );
  AOI21X1 _06365_ (
    .A(clock_module_0.bcsctl2_2_ ),
    .B(_00247_),
    .C(_00248_),
    .Y(_00249_)
  );
  AND2X1 _06366_ (
    .A(_00226_),
    .B(_00249_),
    .Y(_00187_)
  );
  OR2X1 _06367_ (
    .A(clock_module_0.wdt_reset ),
    .B(clock_module_0.por ),
    .Y(clock_module_0.puc_a )
  );
  DFFSR _06368_ (
    .CLK(dco_clk),
    .D(clock_module_0.dbg_rst_nxt ),
    .Q(clock_module_0.dbg_rst ),
    .R(1'h1),
    .S(_00188_)
  );
  DFFSR _06369_ (
    .CLK(dco_clk),
    .D(_00184_),
    .Q(clock_module_0.smclk_div_0_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06370_ (
    .CLK(dco_clk),
    .D(_00185_),
    .Q(clock_module_0.smclk_div_1_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06371_ (
    .CLK(dco_clk),
    .D(_00186_),
    .Q(clock_module_0.smclk_div_2_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06372_ (
    .CLK(dco_clk),
    .D(_00187_),
    .Q(_00163_),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06373_ (
    .CLK(dco_clk),
    .D(_00167_),
    .Q(_00048_),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06374_ (
    .CLK(dco_clk),
    .D(_00164_),
    .Q(clock_module_0.aclk_div_0_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06375_ (
    .CLK(dco_clk),
    .D(_00165_),
    .Q(clock_module_0.aclk_div_1_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06376_ (
    .CLK(dco_clk),
    .D(_00166_),
    .Q(clock_module_0.aclk_div_2_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06377_ (
    .CLK(dco_clk),
    .D(clock_module_0.lfxt_clk_s ),
    .Q(clock_module_0.lfxt_clk_dly ),
    .R(_00188_),
    .S(1'h1)
  );
  DFFSR _06378_ (
    .CLK(dco_clk),
    .D(_00176_),
    .Q(clock_module_0.bcsctl2_0_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06379_ (
    .CLK(dco_clk),
    .D(_00177_),
    .Q(clock_module_0.bcsctl2_1_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06380_ (
    .CLK(dco_clk),
    .D(_00178_),
    .Q(clock_module_0.bcsctl2_2_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06381_ (
    .CLK(dco_clk),
    .D(_00179_),
    .Q(clock_module_0.bcsctl2_3_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06382_ (
    .CLK(dco_clk),
    .D(_00180_),
    .Q(clock_module_0.bcsctl2_4_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06383_ (
    .CLK(dco_clk),
    .D(_00181_),
    .Q(clock_module_0.bcsctl2_5_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06384_ (
    .CLK(dco_clk),
    .D(_00182_),
    .Q(clock_module_0.bcsctl2_6_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06385_ (
    .CLK(dco_clk),
    .D(_00183_),
    .Q(clock_module_0.bcsctl2_7_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06386_ (
    .CLK(dco_clk),
    .D(_00168_),
    .Q(clock_module_0.bcsctl1_0_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06387_ (
    .CLK(dco_clk),
    .D(_00169_),
    .Q(clock_module_0.bcsctl1_1_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06388_ (
    .CLK(dco_clk),
    .D(_00170_),
    .Q(clock_module_0.bcsctl1_2_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06389_ (
    .CLK(dco_clk),
    .D(_00171_),
    .Q(clock_module_0.bcsctl1_3_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06390_ (
    .CLK(dco_clk),
    .D(_00172_),
    .Q(clock_module_0.bcsctl1_4_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06391_ (
    .CLK(dco_clk),
    .D(_00173_),
    .Q(clock_module_0.bcsctl1_5_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06392_ (
    .CLK(dco_clk),
    .D(_00174_),
    .Q(clock_module_0.bcsctl1_6_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  DFFSR _06393_ (
    .CLK(dco_clk),
    .D(_00175_),
    .Q(clock_module_0.bcsctl1_7_ ),
    .R(clock_module_0.puc_noscan_n ),
    .S(1'h1)
  );
  INVX1 _06394_ (
    .A(clock_module_0.por ),
    .Y(_00250_)
  );
  DFFSR _06395_ (
    .CLK(dco_clk),
    .D(lfxt_clk),
    .Q(clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ),
    .R(_00250_),
    .S(1'h1)
  );
  DFFSR _06396_ (
    .CLK(dco_clk),
    .D(clock_module_0.sync_cell_lfxt_clk.data_sync_0_ ),
    .Q(clock_module_0.lfxt_clk_s ),
    .R(_00250_),
    .S(1'h1)
  );
  INVX1 _06397_ (
    .A(clock_module_0.puc_a ),
    .Y(_00251_)
  );
  DFFSR _06398_ (
    .CLK(dco_clk),
    .D(clock_module_0.sync_cell_puc.data_in ),
    .Q(clock_module_0.sync_cell_puc.data_sync_0_ ),
    .R(_00251_),
    .S(1'h1)
  );
  DFFSR _06399_ (
    .CLK(dco_clk),
    .D(clock_module_0.sync_cell_puc.data_sync_0_ ),
    .Q(clock_module_0.puc_noscan_n ),
    .R(_00251_),
    .S(1'h1)
  );
  INVX1 _06400_ (
    .A(clock_module_0.por_a ),
    .Y(_00252_)
  );
  DFFSR _06401_ (
    .CLK(dco_clk),
    .D(1'h0),
    .Q(clock_module_0.sync_reset_por.data_sync_0_ ),
    .R(1'h1),
    .S(_00252_)
  );
  DFFSR _06402_ (
    .CLK(dco_clk),
    .D(clock_module_0.sync_reset_por.data_sync_0_ ),
    .Q(clock_module_0.por ),
    .R(1'h1),
    .S(_00252_)
  );
  INVX1 _06403_ (
    .A(dbg_0.mem_cnt_5_ ),
    .Y(_00321_)
  );
  INVX1 _06404_ (
    .A(dbg_0.mem_cnt_14_ ),
    .Y(_00322_)
  );
  INVX1 _06405_ (
    .A(dbg_0.mem_cnt_10_ ),
    .Y(_00323_)
  );
  INVX1 _06406_ (
    .A(dbg_0.mem_cnt_9_ ),
    .Y(_00324_)
  );
  INVX1 _06407_ (
    .A(dbg_0.mem_start ),
    .Y(_00325_)
  );
  INVX1 _06408_ (
    .A(dbg_0.mem_startb ),
    .Y(_00326_)
  );
  INVX1 _06409_ (
    .A(dbg_0.mem_state_0_ ),
    .Y(_00327_)
  );
  INVX1 _06410_ (
    .A(dbg_0.mem_ctl_1_ ),
    .Y(_00328_)
  );
  INVX1 _06411_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .Y(_00329_)
  );
  INVX1 _06412_ (
    .A(dbg_0.dbg_addr_0_ ),
    .Y(_00330_)
  );
  INVX1 _06413_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00331_)
  );
  INVX1 _06414_ (
    .A(dbg_0.dbg_din_2_ ),
    .Y(_00332_)
  );
  INVX1 _06415_ (
    .A(dbg_0.dbg_din_3_ ),
    .Y(_00333_)
  );
  INVX1 _06416_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .Y(_00334_)
  );
  INVX1 _06417_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .Y(_00335_)
  );
  INVX1 _06418_ (
    .A(dbg_0.dbg_mem_rd_dly ),
    .Y(_00336_)
  );
  INVX1 _06419_ (
    .A(dbg_0.mem_data_8_ ),
    .Y(_00337_)
  );
  INVX1 _06420_ (
    .A(dbg_0.mem_data_9_ ),
    .Y(_00338_)
  );
  INVX1 _06421_ (
    .A(dbg_0.mem_data_10_ ),
    .Y(_00339_)
  );
  INVX1 _06422_ (
    .A(dbg_0.mem_data_11_ ),
    .Y(_00340_)
  );
  INVX1 _06423_ (
    .A(dbg_0.mem_data_12_ ),
    .Y(_00341_)
  );
  INVX1 _06424_ (
    .A(dbg_0.mem_data_13_ ),
    .Y(_00342_)
  );
  INVX1 _06425_ (
    .A(dbg_0.mem_data_14_ ),
    .Y(_00343_)
  );
  INVX1 _06426_ (
    .A(dbg_0.mem_data_15_ ),
    .Y(_00344_)
  );
  INVX1 _06427_ (
    .A(dbg_0.dbg_din_15_ ),
    .Y(_00345_)
  );
  INVX1 _06428_ (
    .A(dbg_0.dbg_rd_rdy ),
    .Y(_00346_)
  );
  INVX1 _06429_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .Y(_00347_)
  );
  INVX1 _06430_ (
    .A(dbg_0.dbg_mem_addr_2_ ),
    .Y(_00348_)
  );
  INVX1 _06431_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .Y(_00349_)
  );
  INVX1 _06432_ (
    .A(dbg_0.dbg_mem_addr_4_ ),
    .Y(_00350_)
  );
  INVX1 _06433_ (
    .A(dbg_0.dbg_mem_addr_7_ ),
    .Y(_00351_)
  );
  INVX1 _06434_ (
    .A(dbg_0.dbg_mem_addr_8_ ),
    .Y(_00352_)
  );
  INVX1 _06435_ (
    .A(dbg_0.dbg_mem_addr_11_ ),
    .Y(_00353_)
  );
  INVX1 _06436_ (
    .A(dbg_0.dbg_mem_addr_12_ ),
    .Y(_00354_)
  );
  INVX1 _06437_ (
    .A(cpu_en),
    .Y(_00355_)
  );
  INVX1 _06438_ (
    .A(clock_module_0.dbg_rst ),
    .Y(_00320_)
  );
  NOR2X1 _06439_ (
    .A(dbg_0.mem_cnt_4_ ),
    .B(dbg_0.mem_cnt_5_ ),
    .Y(_00356_)
  );
  NOR2X1 _06440_ (
    .A(dbg_0.mem_cnt_6_ ),
    .B(dbg_0.mem_cnt_7_ ),
    .Y(_00357_)
  );
  AND2X1 _06441_ (
    .A(_00356_),
    .B(_00357_),
    .Y(_00358_)
  );
  OR2X1 _06442_ (
    .A(dbg_0.mem_cnt_14_ ),
    .B(dbg_0.mem_cnt_15_ ),
    .Y(_00359_)
  );
  OR2X1 _06443_ (
    .A(dbg_0.mem_cnt_12_ ),
    .B(dbg_0.mem_cnt_13_ ),
    .Y(_00360_)
  );
  OR2X1 _06444_ (
    .A(dbg_0.mem_cnt_8_ ),
    .B(dbg_0.mem_cnt_9_ ),
    .Y(_00361_)
  );
  OR2X1 _06445_ (
    .A(dbg_0.mem_cnt_10_ ),
    .B(dbg_0.mem_cnt_11_ ),
    .Y(_00362_)
  );
  OR2X1 _06446_ (
    .A(_00361_),
    .B(_00362_),
    .Y(_00363_)
  );
  OR2X1 _06447_ (
    .A(dbg_0.mem_cnt_3_ ),
    .B(dbg_0.mem_cnt_0_ ),
    .Y(_00364_)
  );
  OR2X1 _06448_ (
    .A(dbg_0.mem_cnt_2_ ),
    .B(dbg_0.mem_cnt_1_ ),
    .Y(_00365_)
  );
  NOR2X1 _06449_ (
    .A(_00364_),
    .B(_00365_),
    .Y(_00366_)
  );
  NOR3X1 _06450_ (
    .A(_00359_),
    .B(_00361_),
    .C(_00362_),
    .Y(_00367_)
  );
  NOR3X1 _06451_ (
    .A(_00360_),
    .B(_00364_),
    .C(_00365_),
    .Y(_00368_)
  );
  NAND3X1 _06452_ (
    .A(_00358_),
    .B(_00367_),
    .C(_00368_),
    .Y(_00369_)
  );
  OAI21X1 _06453_ (
    .A(_00325_),
    .B(_00369_),
    .C(_00326_),
    .Y(_00370_)
  );
  AND2X1 _06454_ (
    .A(dbg_0.mem_state_0_ ),
    .B(_00370_),
    .Y(_00371_)
  );
  AND2X1 _06455_ (
    .A(cpu_halt_st),
    .B(_00371_),
    .Y(_00317_)
  );
  AND2X1 _06456_ (
    .A(cpu_halt_st),
    .B(dbg_0.mem_state_2_ ),
    .Y(_00316_)
  );
  NOR2X1 _06457_ (
    .A(dbg_0.mem_state_2_ ),
    .B(_00371_),
    .Y(_00372_)
  );
  NOR2X1 _06458_ (
    .A(cpu_halt_st),
    .B(_00372_),
    .Y(_00319_)
  );
  NOR2X1 _06459_ (
    .A(dbg_0.mem_state_1_ ),
    .B(dbg_0.mem_state_3_ ),
    .Y(_00373_)
  );
  OAI21X1 _06460_ (
    .A(_00327_),
    .B(_00370_),
    .C(_00373_),
    .Y(_00318_)
  );
  NOR2X1 _06461_ (
    .A(dbg_0.mem_ctl_2_ ),
    .B(_00373_),
    .Y(dbg_0.dbg_mem_en )
  );
  OAI21X1 _06462_ (
    .A(dbg_0.mem_state_1_ ),
    .B(dbg_0.mem_state_3_ ),
    .C(dbg_0.mem_ctl_1_ ),
    .Y(_00374_)
  );
  NAND2X1 _06463_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(dbg_0.dbg_mem_en ),
    .Y(_00375_)
  );
  AOI21X1 _06464_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00329_),
    .C(_00375_),
    .Y(dbg_0.dbg_mem_wr_1_ )
  );
  AND2X1 _06465_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(dbg_0.dbg_mem_addr_0_ ),
    .Y(_00376_)
  );
  NAND2X1 _06466_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(dbg_0.dbg_mem_addr_0_ ),
    .Y(_00377_)
  );
  NOR2X1 _06467_ (
    .A(_00375_),
    .B(_00376_),
    .Y(dbg_0.dbg_mem_wr_0_ )
  );
  OR2X1 _06468_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_addr_1_ ),
    .Y(_00378_)
  );
  OR2X1 _06469_ (
    .A(dbg_0.dbg_addr_0_ ),
    .B(_00378_),
    .Y(_00379_)
  );
  OR2X1 _06470_ (
    .A(dbg_0.dbg_addr_3_ ),
    .B(dbg_0.dbg_addr_4_ ),
    .Y(_00380_)
  );
  NOR2X1 _06471_ (
    .A(dbg_0.dbg_addr_5_ ),
    .B(_00380_),
    .Y(_00381_)
  );
  NAND2X1 _06472_ (
    .A(dbg_0.dbg_addr_2_ ),
    .B(_00381_),
    .Y(_00382_)
  );
  NOR2X1 _06473_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_addr_2_ ),
    .Y(_00383_)
  );
  NOR2X1 _06474_ (
    .A(_00379_),
    .B(_00382_),
    .Y(_00384_)
  );
  AND2X1 _06475_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00384_),
    .Y(_00385_)
  );
  MUX2X1 _06476_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(dbg_0.mem_ctl_1_ ),
    .S(_00385_),
    .Y(_00386_)
  );
  INVX1 _06477_ (
    .A(_00386_),
    .Y(_00295_)
  );
  NAND2X1 _06478_ (
    .A(_00332_),
    .B(_00385_),
    .Y(_00387_)
  );
  OAI21X1 _06479_ (
    .A(dbg_0.mem_ctl_2_ ),
    .B(_00385_),
    .C(_00387_),
    .Y(_00388_)
  );
  INVX1 _06480_ (
    .A(_00388_),
    .Y(_00296_)
  );
  NAND2X1 _06481_ (
    .A(_00333_),
    .B(_00385_),
    .Y(_00389_)
  );
  OAI21X1 _06482_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00385_),
    .C(_00389_),
    .Y(_00390_)
  );
  INVX1 _06483_ (
    .A(_00390_),
    .Y(_00297_)
  );
  NAND3X1 _06484_ (
    .A(dbg_0.dbg_addr_0_ ),
    .B(_00331_),
    .C(dbg_0.dbg_addr_1_ ),
    .Y(_00391_)
  );
  NAND2X1 _06485_ (
    .A(_00381_),
    .B(_00383_),
    .Y(_00392_)
  );
  NOR2X1 _06486_ (
    .A(_00391_),
    .B(_00392_),
    .Y(_00393_)
  );
  NAND2X1 _06487_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00393_),
    .Y(_00394_)
  );
  OR2X1 _06488_ (
    .A(_00332_),
    .B(_00394_),
    .Y(_00395_)
  );
  AOI21X1 _06489_ (
    .A(dbg_0.cpu_stat_2_ ),
    .B(_00395_),
    .C(_00162_),
    .Y(_00396_)
  );
  INVX1 _06490_ (
    .A(_00396_),
    .Y(_00257_)
  );
  OAI21X1 _06491_ (
    .A(_00333_),
    .B(_00394_),
    .C(dbg_0.cpu_stat_3_ ),
    .Y(_00397_)
  );
  NOR2X1 _06492_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .B(dbg_0.fe_mdb_in_5_ ),
    .Y(_00398_)
  );
  NOR2X1 _06493_ (
    .A(dbg_0.fe_mdb_in_3_ ),
    .B(dbg_0.fe_mdb_in_4_ ),
    .Y(_00399_)
  );
  NAND3X1 _06494_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(dbg_0.fe_mdb_in_0_ ),
    .C(_00399_),
    .Y(_00400_)
  );
  INVX1 _06495_ (
    .A(_00400_),
    .Y(_00401_)
  );
  NOR2X1 _06496_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_00335_),
    .Y(_00402_)
  );
  NAND3X1 _06497_ (
    .A(dbg_0.decode_noirq ),
    .B(dbg_0.cpu_ctl_3_ ),
    .C(_00402_),
    .Y(_00403_)
  );
  NOR2X1 _06498_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(dbg_0.fe_mdb_in_12_ ),
    .Y(_00404_)
  );
  NOR2X1 _06499_ (
    .A(dbg_0.fe_mdb_in_11_ ),
    .B(dbg_0.fe_mdb_in_10_ ),
    .Y(_00405_)
  );
  NAND2X1 _06500_ (
    .A(_00334_),
    .B(dbg_0.fe_mdb_in_6_ ),
    .Y(_00406_)
  );
  NAND2X1 _06501_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(dbg_0.fe_mdb_in_8_ ),
    .Y(_00407_)
  );
  NOR2X1 _06502_ (
    .A(_00406_),
    .B(_00407_),
    .Y(_00408_)
  );
  NAND3X1 _06503_ (
    .A(_00404_),
    .B(_00405_),
    .C(_00408_),
    .Y(_00409_)
  );
  NOR2X1 _06504_ (
    .A(_00403_),
    .B(_00409_),
    .Y(_00410_)
  );
  NAND3X1 _06505_ (
    .A(_00398_),
    .B(_00401_),
    .C(_00410_),
    .Y(_00411_)
  );
  NAND2X1 _06506_ (
    .A(_00397_),
    .B(_00411_),
    .Y(_00258_)
  );
  OAI21X1 _06507_ (
    .A(_00330_),
    .B(dbg_0.dbg_i2c_0.mem_burst ),
    .C(_00378_),
    .Y(_00412_)
  );
  NOR2X1 _06508_ (
    .A(_00392_),
    .B(_00412_),
    .Y(_00413_)
  );
  AND2X1 _06509_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00413_),
    .Y(_00414_)
  );
  MUX2X1 _06510_ (
    .A(dbg_0.dbg_din_3_ ),
    .B(dbg_0.cpu_ctl_3_ ),
    .S(_00414_),
    .Y(_00415_)
  );
  INVX1 _06511_ (
    .A(_00415_),
    .Y(_00253_)
  );
  MUX2X1 _06512_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(dbg_0.cpu_ctl_4_ ),
    .S(_00414_),
    .Y(_00416_)
  );
  INVX1 _06513_ (
    .A(_00416_),
    .Y(_00254_)
  );
  MUX2X1 _06514_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(dbg_0.cpu_ctl_5_ ),
    .S(_00414_),
    .Y(_00417_)
  );
  INVX1 _06515_ (
    .A(_00417_),
    .Y(_00255_)
  );
  MUX2X1 _06516_ (
    .A(dbg_0.dbg_din_6_ ),
    .B(clock_module_0.dbg_cpu_reset ),
    .S(_00414_),
    .Y(_00418_)
  );
  INVX1 _06517_ (
    .A(_00418_),
    .Y(_00256_)
  );
  AOI21X1 _06518_ (
    .A(_00331_),
    .B(_00382_),
    .C(_00412_),
    .Y(_00419_)
  );
  AND2X1 _06519_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00419_),
    .Y(_00420_)
  );
  NAND2X1 _06520_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00419_),
    .Y(_00421_)
  );
  OAI21X1 _06521_ (
    .A(dbg_0.mem_state_1_ ),
    .B(dbg_0.mem_state_3_ ),
    .C(dbg_0.mem_ctl_2_ ),
    .Y(_00422_)
  );
  NOR2X1 _06522_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00422_),
    .Y(_00423_)
  );
  NOR2X1 _06523_ (
    .A(dbg_0.dbg_mem_rd_dly ),
    .B(_00423_),
    .Y(_00424_)
  );
  OAI21X1 _06524_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00422_),
    .C(dbg_0.dbg_mem_rd_dly ),
    .Y(_00425_)
  );
  MUX2X1 _06525_ (
    .A(dbg_0.dbg_mem_din_0_ ),
    .B(dbg_0.dbg_mem_din_8_ ),
    .S(_00377_),
    .Y(_00426_)
  );
  NAND2X1 _06526_ (
    .A(dbg_0.dbg_reg_din_0_ ),
    .B(_00423_),
    .Y(_00427_)
  );
  OAI21X1 _06527_ (
    .A(_00425_),
    .B(_00426_),
    .C(_00427_),
    .Y(_00428_)
  );
  AOI21X1 _06528_ (
    .A(dbg_0.mem_data_0_ ),
    .B(_00424_),
    .C(_00428_),
    .Y(_00429_)
  );
  NAND2X1 _06529_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(_00420_),
    .Y(_00430_)
  );
  OAI21X1 _06530_ (
    .A(_00420_),
    .B(_00429_),
    .C(_00430_),
    .Y(_00298_)
  );
  MUX2X1 _06531_ (
    .A(dbg_0.dbg_mem_din_1_ ),
    .B(dbg_0.dbg_mem_din_9_ ),
    .S(_00377_),
    .Y(_00431_)
  );
  NAND2X1 _06532_ (
    .A(dbg_0.dbg_reg_din_1_ ),
    .B(_00423_),
    .Y(_00432_)
  );
  OAI21X1 _06533_ (
    .A(_00425_),
    .B(_00431_),
    .C(_00432_),
    .Y(_00433_)
  );
  AOI21X1 _06534_ (
    .A(dbg_0.mem_data_1_ ),
    .B(_00424_),
    .C(_00433_),
    .Y(_00434_)
  );
  NAND2X1 _06535_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(_00420_),
    .Y(_00435_)
  );
  OAI21X1 _06536_ (
    .A(_00420_),
    .B(_00434_),
    .C(_00435_),
    .Y(_00305_)
  );
  NAND2X1 _06537_ (
    .A(dbg_0.mem_data_2_ ),
    .B(_00424_),
    .Y(_00436_)
  );
  MUX2X1 _06538_ (
    .A(dbg_0.dbg_mem_din_2_ ),
    .B(dbg_0.dbg_mem_din_10_ ),
    .S(_00377_),
    .Y(_00437_)
  );
  AND2X1 _06539_ (
    .A(dbg_0.dbg_reg_din_2_ ),
    .B(_00423_),
    .Y(_00438_)
  );
  OAI21X1 _06540_ (
    .A(_00425_),
    .B(_00437_),
    .C(_00436_),
    .Y(_00439_)
  );
  OAI21X1 _06541_ (
    .A(_00438_),
    .B(_00439_),
    .C(_00421_),
    .Y(_00440_)
  );
  OAI21X1 _06542_ (
    .A(_00332_),
    .B(_00421_),
    .C(_00440_),
    .Y(_00306_)
  );
  NAND2X1 _06543_ (
    .A(dbg_0.mem_data_3_ ),
    .B(_00424_),
    .Y(_00441_)
  );
  MUX2X1 _06544_ (
    .A(dbg_0.dbg_mem_din_3_ ),
    .B(dbg_0.dbg_mem_din_11_ ),
    .S(_00377_),
    .Y(_00442_)
  );
  AND2X1 _06545_ (
    .A(dbg_0.dbg_reg_din_3_ ),
    .B(_00423_),
    .Y(_00443_)
  );
  OAI21X1 _06546_ (
    .A(_00425_),
    .B(_00442_),
    .C(_00441_),
    .Y(_00444_)
  );
  OAI21X1 _06547_ (
    .A(_00443_),
    .B(_00444_),
    .C(_00421_),
    .Y(_00445_)
  );
  OAI21X1 _06548_ (
    .A(_00333_),
    .B(_00421_),
    .C(_00445_),
    .Y(_00307_)
  );
  MUX2X1 _06549_ (
    .A(dbg_0.dbg_mem_din_4_ ),
    .B(dbg_0.dbg_mem_din_12_ ),
    .S(_00377_),
    .Y(_00446_)
  );
  NAND2X1 _06550_ (
    .A(dbg_0.dbg_reg_din_4_ ),
    .B(_00423_),
    .Y(_00447_)
  );
  OAI21X1 _06551_ (
    .A(_00425_),
    .B(_00446_),
    .C(_00447_),
    .Y(_00448_)
  );
  AOI21X1 _06552_ (
    .A(dbg_0.mem_data_4_ ),
    .B(_00424_),
    .C(_00448_),
    .Y(_00449_)
  );
  NAND2X1 _06553_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(_00420_),
    .Y(_00450_)
  );
  OAI21X1 _06554_ (
    .A(_00420_),
    .B(_00449_),
    .C(_00450_),
    .Y(_00308_)
  );
  NAND2X1 _06555_ (
    .A(dbg_0.dbg_reg_din_5_ ),
    .B(_00423_),
    .Y(_00451_)
  );
  MUX2X1 _06556_ (
    .A(dbg_0.dbg_mem_din_5_ ),
    .B(dbg_0.dbg_mem_din_13_ ),
    .S(_00377_),
    .Y(_00452_)
  );
  OAI21X1 _06557_ (
    .A(_00425_),
    .B(_00452_),
    .C(_00451_),
    .Y(_00453_)
  );
  AOI21X1 _06558_ (
    .A(dbg_0.mem_data_5_ ),
    .B(_00424_),
    .C(_00453_),
    .Y(_00454_)
  );
  NAND2X1 _06559_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(_00420_),
    .Y(_00455_)
  );
  OAI21X1 _06560_ (
    .A(_00420_),
    .B(_00454_),
    .C(_00455_),
    .Y(_00309_)
  );
  NAND2X1 _06561_ (
    .A(dbg_0.dbg_reg_din_6_ ),
    .B(_00423_),
    .Y(_00456_)
  );
  MUX2X1 _06562_ (
    .A(dbg_0.dbg_mem_din_6_ ),
    .B(dbg_0.dbg_mem_din_14_ ),
    .S(_00377_),
    .Y(_00457_)
  );
  OAI21X1 _06563_ (
    .A(_00425_),
    .B(_00457_),
    .C(_00456_),
    .Y(_00458_)
  );
  AOI21X1 _06564_ (
    .A(dbg_0.mem_data_6_ ),
    .B(_00424_),
    .C(_00458_),
    .Y(_00459_)
  );
  NAND2X1 _06565_ (
    .A(dbg_0.dbg_din_6_ ),
    .B(_00420_),
    .Y(_00460_)
  );
  OAI21X1 _06566_ (
    .A(_00420_),
    .B(_00459_),
    .C(_00460_),
    .Y(_00310_)
  );
  MUX2X1 _06567_ (
    .A(dbg_0.dbg_mem_din_7_ ),
    .B(dbg_0.dbg_mem_din_15_ ),
    .S(_00377_),
    .Y(_00461_)
  );
  NAND2X1 _06568_ (
    .A(dbg_0.dbg_reg_din_7_ ),
    .B(_00423_),
    .Y(_00462_)
  );
  OAI21X1 _06569_ (
    .A(_00425_),
    .B(_00461_),
    .C(_00462_),
    .Y(_00463_)
  );
  AOI21X1 _06570_ (
    .A(dbg_0.mem_data_7_ ),
    .B(_00424_),
    .C(_00463_),
    .Y(_00464_)
  );
  NAND2X1 _06571_ (
    .A(dbg_0.dbg_din_7_ ),
    .B(_00420_),
    .Y(_00465_)
  );
  OAI21X1 _06572_ (
    .A(_00420_),
    .B(_00464_),
    .C(_00465_),
    .Y(_00311_)
  );
  NOR2X1 _06573_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00336_),
    .Y(_00466_)
  );
  NAND2X1 _06574_ (
    .A(dbg_0.dbg_mem_din_8_ ),
    .B(_00466_),
    .Y(_00467_)
  );
  NAND2X1 _06575_ (
    .A(dbg_0.dbg_reg_din_8_ ),
    .B(_00423_),
    .Y(_00468_)
  );
  OAI21X1 _06576_ (
    .A(_00423_),
    .B(_00467_),
    .C(_00468_),
    .Y(_00469_)
  );
  AOI21X1 _06577_ (
    .A(dbg_0.mem_data_8_ ),
    .B(_00424_),
    .C(_00469_),
    .Y(_00470_)
  );
  NOR2X1 _06578_ (
    .A(dbg_0.dbg_din_8_ ),
    .B(_00421_),
    .Y(_00471_)
  );
  AOI21X1 _06579_ (
    .A(_00421_),
    .B(_00470_),
    .C(_00471_),
    .Y(_00312_)
  );
  NAND2X1 _06580_ (
    .A(dbg_0.dbg_mem_din_9_ ),
    .B(_00466_),
    .Y(_00472_)
  );
  NAND2X1 _06581_ (
    .A(dbg_0.dbg_reg_din_9_ ),
    .B(_00423_),
    .Y(_00473_)
  );
  OAI21X1 _06582_ (
    .A(_00423_),
    .B(_00472_),
    .C(_00473_),
    .Y(_00474_)
  );
  AOI21X1 _06583_ (
    .A(dbg_0.mem_data_9_ ),
    .B(_00424_),
    .C(_00474_),
    .Y(_00475_)
  );
  NOR2X1 _06584_ (
    .A(dbg_0.dbg_din_9_ ),
    .B(_00421_),
    .Y(_00476_)
  );
  AOI21X1 _06585_ (
    .A(_00421_),
    .B(_00475_),
    .C(_00476_),
    .Y(_00313_)
  );
  NAND2X1 _06586_ (
    .A(dbg_0.dbg_mem_din_10_ ),
    .B(_00466_),
    .Y(_00477_)
  );
  NAND2X1 _06587_ (
    .A(dbg_0.dbg_reg_din_10_ ),
    .B(_00423_),
    .Y(_00478_)
  );
  OAI21X1 _06588_ (
    .A(_00423_),
    .B(_00477_),
    .C(_00478_),
    .Y(_00479_)
  );
  AOI21X1 _06589_ (
    .A(dbg_0.mem_data_10_ ),
    .B(_00424_),
    .C(_00479_),
    .Y(_00480_)
  );
  NOR2X1 _06590_ (
    .A(dbg_0.dbg_din_10_ ),
    .B(_00421_),
    .Y(_00481_)
  );
  AOI21X1 _06591_ (
    .A(_00421_),
    .B(_00480_),
    .C(_00481_),
    .Y(_00299_)
  );
  NAND2X1 _06592_ (
    .A(dbg_0.dbg_mem_din_11_ ),
    .B(_00466_),
    .Y(_00482_)
  );
  NAND2X1 _06593_ (
    .A(dbg_0.dbg_reg_din_11_ ),
    .B(_00423_),
    .Y(_00483_)
  );
  OAI21X1 _06594_ (
    .A(_00423_),
    .B(_00482_),
    .C(_00483_),
    .Y(_00484_)
  );
  AOI21X1 _06595_ (
    .A(dbg_0.mem_data_11_ ),
    .B(_00424_),
    .C(_00484_),
    .Y(_00485_)
  );
  NOR2X1 _06596_ (
    .A(dbg_0.dbg_din_11_ ),
    .B(_00421_),
    .Y(_00486_)
  );
  AOI21X1 _06597_ (
    .A(_00421_),
    .B(_00485_),
    .C(_00486_),
    .Y(_00300_)
  );
  NAND2X1 _06598_ (
    .A(dbg_0.dbg_mem_din_12_ ),
    .B(_00466_),
    .Y(_00487_)
  );
  NAND2X1 _06599_ (
    .A(dbg_0.dbg_reg_din_12_ ),
    .B(_00423_),
    .Y(_00488_)
  );
  OAI21X1 _06600_ (
    .A(_00423_),
    .B(_00487_),
    .C(_00488_),
    .Y(_00489_)
  );
  AOI21X1 _06601_ (
    .A(dbg_0.mem_data_12_ ),
    .B(_00424_),
    .C(_00489_),
    .Y(_00490_)
  );
  NOR2X1 _06602_ (
    .A(dbg_0.dbg_din_12_ ),
    .B(_00421_),
    .Y(_00491_)
  );
  AOI21X1 _06603_ (
    .A(_00421_),
    .B(_00490_),
    .C(_00491_),
    .Y(_00301_)
  );
  NAND2X1 _06604_ (
    .A(dbg_0.dbg_mem_din_13_ ),
    .B(_00466_),
    .Y(_00492_)
  );
  NAND2X1 _06605_ (
    .A(dbg_0.dbg_reg_din_13_ ),
    .B(_00423_),
    .Y(_00493_)
  );
  OAI21X1 _06606_ (
    .A(_00423_),
    .B(_00492_),
    .C(_00493_),
    .Y(_00494_)
  );
  AOI21X1 _06607_ (
    .A(dbg_0.mem_data_13_ ),
    .B(_00424_),
    .C(_00494_),
    .Y(_00495_)
  );
  NOR2X1 _06608_ (
    .A(dbg_0.dbg_din_13_ ),
    .B(_00421_),
    .Y(_00496_)
  );
  AOI21X1 _06609_ (
    .A(_00421_),
    .B(_00495_),
    .C(_00496_),
    .Y(_00302_)
  );
  NAND2X1 _06610_ (
    .A(dbg_0.dbg_mem_din_14_ ),
    .B(_00466_),
    .Y(_00497_)
  );
  NAND2X1 _06611_ (
    .A(dbg_0.dbg_reg_din_14_ ),
    .B(_00423_),
    .Y(_00498_)
  );
  OAI21X1 _06612_ (
    .A(_00423_),
    .B(_00497_),
    .C(_00498_),
    .Y(_00499_)
  );
  AOI21X1 _06613_ (
    .A(dbg_0.mem_data_14_ ),
    .B(_00424_),
    .C(_00499_),
    .Y(_00500_)
  );
  NOR2X1 _06614_ (
    .A(dbg_0.dbg_din_14_ ),
    .B(_00421_),
    .Y(_00501_)
  );
  AOI21X1 _06615_ (
    .A(_00421_),
    .B(_00500_),
    .C(_00501_),
    .Y(_00303_)
  );
  NAND2X1 _06616_ (
    .A(dbg_0.dbg_mem_din_15_ ),
    .B(_00466_),
    .Y(_00502_)
  );
  NAND2X1 _06617_ (
    .A(dbg_0.dbg_reg_din_15_ ),
    .B(_00423_),
    .Y(_00503_)
  );
  OAI21X1 _06618_ (
    .A(_00423_),
    .B(_00502_),
    .C(_00503_),
    .Y(_00504_)
  );
  AOI21X1 _06619_ (
    .A(dbg_0.mem_data_15_ ),
    .B(_00424_),
    .C(_00504_),
    .Y(_00505_)
  );
  MUX2X1 _06620_ (
    .A(_00345_),
    .B(_00505_),
    .S(_00420_),
    .Y(_00304_)
  );
  NAND2X1 _06621_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(_00414_),
    .Y(_00506_)
  );
  AND2X1 _06622_ (
    .A(dbg_0.cpu_ctl_5_ ),
    .B(dbg_en),
    .Y(_00507_)
  );
  AOI21X1 _06623_ (
    .A(_00162_),
    .B(_00507_),
    .C(dbg_0.halt_flag ),
    .Y(_00508_)
  );
  AND2X1 _06624_ (
    .A(_00411_),
    .B(_00508_),
    .Y(_00509_)
  );
  OAI21X1 _06625_ (
    .A(cpu_halt_st),
    .B(_00506_),
    .C(_00509_),
    .Y(_00510_)
  );
  AOI21X1 _06626_ (
    .A(dbg_0.mem_state_0_ ),
    .B(_00319_),
    .C(_00510_),
    .Y(_00511_)
  );
  NAND3X1 _06627_ (
    .A(cpu_halt_st),
    .B(dbg_0.dbg_din_1_ ),
    .C(_00414_),
    .Y(_00512_)
  );
  AOI21X1 _06628_ (
    .A(dbg_0.mem_state_1_ ),
    .B(_00372_),
    .C(_00511_),
    .Y(_00513_)
  );
  AND2X1 _06629_ (
    .A(_00512_),
    .B(_00513_),
    .Y(_00260_)
  );
  OR2X1 _06630_ (
    .A(_00330_),
    .B(_00378_),
    .Y(_00514_)
  );
  NOR2X1 _06631_ (
    .A(_00382_),
    .B(_00514_),
    .Y(_00515_)
  );
  AND2X1 _06632_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00515_),
    .Y(_00516_)
  );
  NAND2X1 _06633_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00515_),
    .Y(_00517_)
  );
  AOI21X1 _06634_ (
    .A(_00346_),
    .B(_00374_),
    .C(_00331_),
    .Y(_00518_)
  );
  AND2X1 _06635_ (
    .A(_00369_),
    .B(_00518_),
    .Y(_00519_)
  );
  NAND2X1 _06636_ (
    .A(_00369_),
    .B(_00518_),
    .Y(_00520_)
  );
  OR2X1 _06637_ (
    .A(dbg_0.mem_ctl_2_ ),
    .B(dbg_0.dbg_i2c_0.mem_bw ),
    .Y(_00521_)
  );
  NAND3X1 _06638_ (
    .A(_00369_),
    .B(_00518_),
    .C(_00521_),
    .Y(_00522_)
  );
  OR2X1 _06639_ (
    .A(_00329_),
    .B(_00522_),
    .Y(_00523_)
  );
  NAND2X1 _06640_ (
    .A(_00329_),
    .B(_00522_),
    .Y(_00524_)
  );
  NAND2X1 _06641_ (
    .A(_00523_),
    .B(_00524_),
    .Y(_00525_)
  );
  NAND2X1 _06642_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(_00516_),
    .Y(_00526_)
  );
  OAI21X1 _06643_ (
    .A(_00516_),
    .B(_00525_),
    .C(_00526_),
    .Y(_00262_)
  );
  NOR2X1 _06644_ (
    .A(_00520_),
    .B(_00521_),
    .Y(_00527_)
  );
  NOR3X1 _06645_ (
    .A(_00347_),
    .B(_00520_),
    .C(_00521_),
    .Y(_00528_)
  );
  NOR2X1 _06646_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .B(_00527_),
    .Y(_00529_)
  );
  OAI21X1 _06647_ (
    .A(_00528_),
    .B(_00529_),
    .C(_00523_),
    .Y(_00530_)
  );
  NOR3X1 _06648_ (
    .A(_00329_),
    .B(_00347_),
    .C(_00522_),
    .Y(_00531_)
  );
  OAI21X1 _06649_ (
    .A(_00347_),
    .B(_00523_),
    .C(_00530_),
    .Y(_00532_)
  );
  NAND2X1 _06650_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(_00516_),
    .Y(_00533_)
  );
  OAI21X1 _06651_ (
    .A(_00516_),
    .B(_00532_),
    .C(_00533_),
    .Y(_00269_)
  );
  NOR2X1 _06652_ (
    .A(_00528_),
    .B(_00531_),
    .Y(_00534_)
  );
  OAI21X1 _06653_ (
    .A(_00528_),
    .B(_00531_),
    .C(dbg_0.dbg_mem_addr_2_ ),
    .Y(_00535_)
  );
  NAND2X1 _06654_ (
    .A(_00348_),
    .B(_00534_),
    .Y(_00536_)
  );
  AOI21X1 _06655_ (
    .A(_00535_),
    .B(_00536_),
    .C(_00516_),
    .Y(_00537_)
  );
  AOI21X1 _06656_ (
    .A(_00332_),
    .B(_00516_),
    .C(_00537_),
    .Y(_00270_)
  );
  XNOR2X1 _06657_ (
    .A(_00349_),
    .B(_00535_),
    .Y(_00538_)
  );
  MUX2X1 _06658_ (
    .A(_00333_),
    .B(_00538_),
    .S(_00516_),
    .Y(_00271_)
  );
  OAI21X1 _06659_ (
    .A(_00349_),
    .B(_00535_),
    .C(_00350_),
    .Y(_00539_)
  );
  INVX1 _06660_ (
    .A(_00539_),
    .Y(_00540_)
  );
  NOR3X1 _06661_ (
    .A(_00349_),
    .B(_00350_),
    .C(_00535_),
    .Y(_00541_)
  );
  OR2X1 _06662_ (
    .A(_00540_),
    .B(_00541_),
    .Y(_00542_)
  );
  NAND2X1 _06663_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(_00516_),
    .Y(_00543_)
  );
  OAI21X1 _06664_ (
    .A(_00516_),
    .B(_00542_),
    .C(_00543_),
    .Y(_00272_)
  );
  NAND2X1 _06665_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(_00516_),
    .Y(_00544_)
  );
  XNOR2X1 _06666_ (
    .A(dbg_0.dbg_mem_addr_5_ ),
    .B(_00541_),
    .Y(_00545_)
  );
  OAI21X1 _06667_ (
    .A(_00516_),
    .B(_00545_),
    .C(_00544_),
    .Y(_00273_)
  );
  NAND3X1 _06668_ (
    .A(dbg_0.dbg_mem_addr_5_ ),
    .B(dbg_0.dbg_mem_addr_6_ ),
    .C(_00541_),
    .Y(_00546_)
  );
  AOI21X1 _06669_ (
    .A(dbg_0.dbg_mem_addr_5_ ),
    .B(_00541_),
    .C(dbg_0.dbg_mem_addr_6_ ),
    .Y(_00547_)
  );
  INVX1 _06670_ (
    .A(_00547_),
    .Y(_00548_)
  );
  NOR2X1 _06671_ (
    .A(dbg_0.dbg_din_6_ ),
    .B(_00517_),
    .Y(_00549_)
  );
  AOI21X1 _06672_ (
    .A(_00546_),
    .B(_00548_),
    .C(_00516_),
    .Y(_00550_)
  );
  NOR2X1 _06673_ (
    .A(_00549_),
    .B(_00550_),
    .Y(_00274_)
  );
  NAND2X1 _06674_ (
    .A(dbg_0.dbg_din_7_ ),
    .B(_00516_),
    .Y(_00551_)
  );
  XNOR2X1 _06675_ (
    .A(_00351_),
    .B(_00546_),
    .Y(_00552_)
  );
  OAI21X1 _06676_ (
    .A(_00516_),
    .B(_00552_),
    .C(_00551_),
    .Y(_00275_)
  );
  NAND2X1 _06677_ (
    .A(dbg_0.dbg_din_8_ ),
    .B(_00516_),
    .Y(_00553_)
  );
  NOR3X1 _06678_ (
    .A(_00351_),
    .B(_00352_),
    .C(_00546_),
    .Y(_00554_)
  );
  OAI21X1 _06679_ (
    .A(_00351_),
    .B(_00546_),
    .C(_00352_),
    .Y(_00555_)
  );
  NAND2X1 _06680_ (
    .A(_00517_),
    .B(_00555_),
    .Y(_00556_)
  );
  OAI21X1 _06681_ (
    .A(_00554_),
    .B(_00556_),
    .C(_00553_),
    .Y(_00276_)
  );
  NAND2X1 _06682_ (
    .A(dbg_0.dbg_din_9_ ),
    .B(_00516_),
    .Y(_00557_)
  );
  NAND2X1 _06683_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .B(_00554_),
    .Y(_00558_)
  );
  XNOR2X1 _06684_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .B(_00554_),
    .Y(_00559_)
  );
  OAI21X1 _06685_ (
    .A(_00516_),
    .B(_00559_),
    .C(_00557_),
    .Y(_00277_)
  );
  NAND2X1 _06686_ (
    .A(dbg_0.dbg_din_10_ ),
    .B(_00516_),
    .Y(_00560_)
  );
  NAND3X1 _06687_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .B(dbg_0.dbg_mem_addr_10_ ),
    .C(_00554_),
    .Y(_00561_)
  );
  XOR2X1 _06688_ (
    .A(dbg_0.dbg_mem_addr_10_ ),
    .B(_00558_),
    .Y(_00562_)
  );
  OAI21X1 _06689_ (
    .A(_00516_),
    .B(_00562_),
    .C(_00560_),
    .Y(_00263_)
  );
  NAND2X1 _06690_ (
    .A(dbg_0.dbg_din_11_ ),
    .B(_00516_),
    .Y(_00563_)
  );
  XNOR2X1 _06691_ (
    .A(_00353_),
    .B(_00561_),
    .Y(_00564_)
  );
  OAI21X1 _06692_ (
    .A(_00516_),
    .B(_00564_),
    .C(_00563_),
    .Y(_00264_)
  );
  NAND2X1 _06693_ (
    .A(dbg_0.dbg_din_12_ ),
    .B(_00516_),
    .Y(_00565_)
  );
  NOR3X1 _06694_ (
    .A(_00353_),
    .B(_00354_),
    .C(_00561_),
    .Y(_00566_)
  );
  OAI21X1 _06695_ (
    .A(_00353_),
    .B(_00561_),
    .C(_00354_),
    .Y(_00567_)
  );
  NAND2X1 _06696_ (
    .A(_00517_),
    .B(_00567_),
    .Y(_00568_)
  );
  OAI21X1 _06697_ (
    .A(_00566_),
    .B(_00568_),
    .C(_00565_),
    .Y(_00265_)
  );
  NAND2X1 _06698_ (
    .A(dbg_0.dbg_din_13_ ),
    .B(_00516_),
    .Y(_00569_)
  );
  NAND2X1 _06699_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .B(_00566_),
    .Y(_00570_)
  );
  XNOR2X1 _06700_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .B(_00566_),
    .Y(_00571_)
  );
  OAI21X1 _06701_ (
    .A(_00516_),
    .B(_00571_),
    .C(_00569_),
    .Y(_00266_)
  );
  NAND2X1 _06702_ (
    .A(dbg_0.dbg_din_14_ ),
    .B(_00516_),
    .Y(_00572_)
  );
  NAND3X1 _06703_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .B(dbg_0.dbg_mem_addr_14_ ),
    .C(_00566_),
    .Y(_00573_)
  );
  XOR2X1 _06704_ (
    .A(dbg_0.dbg_mem_addr_14_ ),
    .B(_00570_),
    .Y(_00574_)
  );
  OAI21X1 _06705_ (
    .A(_00516_),
    .B(_00574_),
    .C(_00572_),
    .Y(_00267_)
  );
  OR2X1 _06706_ (
    .A(dbg_0.dbg_mem_addr_15_ ),
    .B(_00573_),
    .Y(_00575_)
  );
  AOI21X1 _06707_ (
    .A(dbg_0.dbg_mem_addr_15_ ),
    .B(_00573_),
    .C(_00516_),
    .Y(_00576_)
  );
  AOI22X1 _06708_ (
    .A(_00345_),
    .B(_00516_),
    .C(_00575_),
    .D(_00576_),
    .Y(_00268_)
  );
  NAND2X1 _06709_ (
    .A(dbg_0.mem_start ),
    .B(_00369_),
    .Y(_00577_)
  );
  NOR2X1 _06710_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00577_),
    .Y(dbg_0.dbg_i2c_0.mem_burst_rd )
  );
  NOR2X1 _06711_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_i2c_0.mem_burst_rd ),
    .Y(_00578_)
  );
  NAND2X1 _06712_ (
    .A(dbg_0.dbg_i2c_0.dbg_rd ),
    .B(_00578_),
    .Y(_00579_)
  );
  OAI21X1 _06713_ (
    .A(_00424_),
    .B(_00578_),
    .C(_00579_),
    .Y(_00259_)
  );
  NAND3X1 _06714_ (
    .A(cpu_halt_st),
    .B(dbg_0.dbg_din_2_ ),
    .C(_00414_),
    .Y(_00580_)
  );
  INVX1 _06715_ (
    .A(_00580_),
    .Y(dbg_0.istep )
  );
  OR2X1 _06716_ (
    .A(dbg_0.inc_step_0_ ),
    .B(dbg_0.istep ),
    .Y(_00261_)
  );
  NOR2X1 _06717_ (
    .A(_00382_),
    .B(_00391_),
    .Y(_00581_)
  );
  AND2X1 _06718_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00581_),
    .Y(_00582_)
  );
  NAND2X1 _06719_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(_00581_),
    .Y(_00583_)
  );
  OR2X1 _06720_ (
    .A(dbg_0.mem_cnt_0_ ),
    .B(_00520_),
    .Y(_00584_)
  );
  XNOR2X1 _06721_ (
    .A(dbg_0.mem_cnt_0_ ),
    .B(_00519_),
    .Y(_00585_)
  );
  NAND2X1 _06722_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(_00582_),
    .Y(_00586_)
  );
  OAI21X1 _06723_ (
    .A(_00582_),
    .B(_00585_),
    .C(_00586_),
    .Y(_00279_)
  );
  NOR2X1 _06724_ (
    .A(dbg_0.mem_cnt_1_ ),
    .B(_00584_),
    .Y(_00587_)
  );
  XOR2X1 _06725_ (
    .A(dbg_0.mem_cnt_1_ ),
    .B(_00584_),
    .Y(_00588_)
  );
  NAND2X1 _06726_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(_00582_),
    .Y(_00589_)
  );
  OAI21X1 _06727_ (
    .A(_00582_),
    .B(_00588_),
    .C(_00589_),
    .Y(_00286_)
  );
  NAND2X1 _06728_ (
    .A(dbg_0.dbg_din_2_ ),
    .B(_00582_),
    .Y(_00590_)
  );
  XNOR2X1 _06729_ (
    .A(dbg_0.mem_cnt_2_ ),
    .B(_00587_),
    .Y(_00591_)
  );
  OAI21X1 _06730_ (
    .A(_00582_),
    .B(_00591_),
    .C(_00590_),
    .Y(_00287_)
  );
  OAI21X1 _06731_ (
    .A(_00365_),
    .B(_00584_),
    .C(dbg_0.mem_cnt_3_ ),
    .Y(_00592_)
  );
  NAND2X1 _06732_ (
    .A(_00366_),
    .B(_00519_),
    .Y(_00593_)
  );
  NAND3X1 _06733_ (
    .A(_00583_),
    .B(_00592_),
    .C(_00593_),
    .Y(_00594_)
  );
  OAI21X1 _06734_ (
    .A(dbg_0.dbg_din_3_ ),
    .B(_00583_),
    .C(_00594_),
    .Y(_00595_)
  );
  INVX1 _06735_ (
    .A(_00595_),
    .Y(_00288_)
  );
  NOR2X1 _06736_ (
    .A(dbg_0.mem_cnt_4_ ),
    .B(_00593_),
    .Y(_00596_)
  );
  XOR2X1 _06737_ (
    .A(dbg_0.mem_cnt_4_ ),
    .B(_00593_),
    .Y(_00597_)
  );
  NAND2X1 _06738_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(_00582_),
    .Y(_00598_)
  );
  OAI21X1 _06739_ (
    .A(_00582_),
    .B(_00597_),
    .C(_00598_),
    .Y(_00289_)
  );
  XNOR2X1 _06740_ (
    .A(dbg_0.mem_cnt_5_ ),
    .B(_00596_),
    .Y(_00599_)
  );
  NAND2X1 _06741_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(_00582_),
    .Y(_00600_)
  );
  OAI21X1 _06742_ (
    .A(_00582_),
    .B(_00599_),
    .C(_00600_),
    .Y(_00290_)
  );
  NAND3X1 _06743_ (
    .A(_00356_),
    .B(_00366_),
    .C(_00519_),
    .Y(_00601_)
  );
  NOR2X1 _06744_ (
    .A(dbg_0.mem_cnt_6_ ),
    .B(_00601_),
    .Y(_00602_)
  );
  XOR2X1 _06745_ (
    .A(dbg_0.mem_cnt_6_ ),
    .B(_00601_),
    .Y(_00603_)
  );
  NAND2X1 _06746_ (
    .A(dbg_0.dbg_din_6_ ),
    .B(_00582_),
    .Y(_00604_)
  );
  OAI21X1 _06747_ (
    .A(_00582_),
    .B(_00603_),
    .C(_00604_),
    .Y(_00291_)
  );
  XNOR2X1 _06748_ (
    .A(dbg_0.mem_cnt_7_ ),
    .B(_00602_),
    .Y(_00605_)
  );
  NAND2X1 _06749_ (
    .A(dbg_0.dbg_din_7_ ),
    .B(_00582_),
    .Y(_00606_)
  );
  OAI21X1 _06750_ (
    .A(_00582_),
    .B(_00605_),
    .C(_00606_),
    .Y(_00292_)
  );
  OR2X1 _06751_ (
    .A(dbg_0.mem_cnt_4_ ),
    .B(_00366_),
    .Y(_00607_)
  );
  AND2X1 _06752_ (
    .A(dbg_0.mem_cnt_6_ ),
    .B(dbg_0.mem_cnt_7_ ),
    .Y(_00608_)
  );
  OAI21X1 _06753_ (
    .A(dbg_0.mem_cnt_7_ ),
    .B(_00520_),
    .C(_00321_),
    .Y(_00609_)
  );
  OAI21X1 _06754_ (
    .A(_00321_),
    .B(_00608_),
    .C(_00609_),
    .Y(_00610_)
  );
  OAI21X1 _06755_ (
    .A(_00607_),
    .B(_00610_),
    .C(_00358_),
    .Y(_00611_)
  );
  OR2X1 _06756_ (
    .A(_00520_),
    .B(_00611_),
    .Y(_00612_)
  );
  NOR2X1 _06757_ (
    .A(dbg_0.mem_cnt_8_ ),
    .B(_00612_),
    .Y(_00613_)
  );
  XOR2X1 _06758_ (
    .A(dbg_0.mem_cnt_8_ ),
    .B(_00612_),
    .Y(_00614_)
  );
  NAND2X1 _06759_ (
    .A(dbg_0.dbg_din_8_ ),
    .B(_00582_),
    .Y(_00615_)
  );
  OAI21X1 _06760_ (
    .A(_00582_),
    .B(_00614_),
    .C(_00615_),
    .Y(_00293_)
  );
  NOR2X1 _06761_ (
    .A(dbg_0.dbg_din_9_ ),
    .B(_00583_),
    .Y(_00616_)
  );
  OAI21X1 _06762_ (
    .A(dbg_0.mem_cnt_8_ ),
    .B(_00612_),
    .C(dbg_0.mem_cnt_9_ ),
    .Y(_00617_)
  );
  NAND2X1 _06763_ (
    .A(_00324_),
    .B(_00613_),
    .Y(_00618_)
  );
  AOI21X1 _06764_ (
    .A(_00324_),
    .B(_00613_),
    .C(_00582_),
    .Y(_00619_)
  );
  AOI21X1 _06765_ (
    .A(_00617_),
    .B(_00619_),
    .C(_00616_),
    .Y(_00294_)
  );
  NAND2X1 _06766_ (
    .A(dbg_0.dbg_din_10_ ),
    .B(_00582_),
    .Y(_00620_)
  );
  NOR2X1 _06767_ (
    .A(dbg_0.mem_cnt_10_ ),
    .B(_00618_),
    .Y(_00621_)
  );
  XNOR2X1 _06768_ (
    .A(_00323_),
    .B(_00618_),
    .Y(_00622_)
  );
  OAI21X1 _06769_ (
    .A(_00582_),
    .B(_00622_),
    .C(_00620_),
    .Y(_00280_)
  );
  NAND2X1 _06770_ (
    .A(dbg_0.dbg_din_11_ ),
    .B(_00582_),
    .Y(_00623_)
  );
  NOR2X1 _06771_ (
    .A(dbg_0.mem_cnt_11_ ),
    .B(_00621_),
    .Y(_00624_)
  );
  OAI21X1 _06772_ (
    .A(_00323_),
    .B(_00520_),
    .C(dbg_0.mem_cnt_11_ ),
    .Y(_00625_)
  );
  OAI21X1 _06773_ (
    .A(_00618_),
    .B(_00625_),
    .C(_00583_),
    .Y(_00626_)
  );
  OAI21X1 _06774_ (
    .A(_00624_),
    .B(_00626_),
    .C(_00623_),
    .Y(_00281_)
  );
  NAND2X1 _06775_ (
    .A(dbg_0.dbg_din_12_ ),
    .B(_00582_),
    .Y(_00627_)
  );
  NAND2X1 _06776_ (
    .A(dbg_0.mem_cnt_12_ ),
    .B(_00519_),
    .Y(_00628_)
  );
  XNOR2X1 _06777_ (
    .A(dbg_0.mem_cnt_12_ ),
    .B(_00519_),
    .Y(_00629_)
  );
  OAI21X1 _06778_ (
    .A(_00363_),
    .B(_00611_),
    .C(_00518_),
    .Y(_00630_)
  );
  XNOR2X1 _06779_ (
    .A(_00629_),
    .B(_00630_),
    .Y(_00631_)
  );
  OAI21X1 _06780_ (
    .A(_00582_),
    .B(_00631_),
    .C(_00627_),
    .Y(_00282_)
  );
  NOR2X1 _06781_ (
    .A(dbg_0.dbg_din_13_ ),
    .B(_00583_),
    .Y(_00632_)
  );
  OAI21X1 _06782_ (
    .A(_00629_),
    .B(_00630_),
    .C(_00628_),
    .Y(_00633_)
  );
  NOR2X1 _06783_ (
    .A(dbg_0.mem_cnt_13_ ),
    .B(_00519_),
    .Y(_00634_)
  );
  AND2X1 _06784_ (
    .A(dbg_0.mem_cnt_13_ ),
    .B(_00519_),
    .Y(_00635_)
  );
  NOR2X1 _06785_ (
    .A(_00634_),
    .B(_00635_),
    .Y(_00636_)
  );
  XNOR2X1 _06786_ (
    .A(_00633_),
    .B(_00636_),
    .Y(_00637_)
  );
  AOI21X1 _06787_ (
    .A(_00583_),
    .B(_00637_),
    .C(_00632_),
    .Y(_00283_)
  );
  NAND2X1 _06788_ (
    .A(dbg_0.dbg_din_14_ ),
    .B(_00582_),
    .Y(_00638_)
  );
  XNOR2X1 _06789_ (
    .A(_00322_),
    .B(_00519_),
    .Y(_00639_)
  );
  NOR2X1 _06790_ (
    .A(_00633_),
    .B(_00635_),
    .Y(_00640_)
  );
  OAI21X1 _06791_ (
    .A(_00633_),
    .B(_00635_),
    .C(_00639_),
    .Y(_00641_)
  );
  XOR2X1 _06792_ (
    .A(_00639_),
    .B(_00640_),
    .Y(_00642_)
  );
  OAI21X1 _06793_ (
    .A(_00582_),
    .B(_00642_),
    .C(_00638_),
    .Y(_00284_)
  );
  OAI21X1 _06794_ (
    .A(_00322_),
    .B(_00520_),
    .C(_00641_),
    .Y(_00643_)
  );
  XNOR2X1 _06795_ (
    .A(dbg_0.mem_cnt_15_ ),
    .B(_00520_),
    .Y(_00644_)
  );
  XNOR2X1 _06796_ (
    .A(_00643_),
    .B(_00644_),
    .Y(_00645_)
  );
  NAND2X1 _06797_ (
    .A(dbg_0.dbg_din_15_ ),
    .B(_00582_),
    .Y(_00646_)
  );
  OAI21X1 _06798_ (
    .A(_00582_),
    .B(_00645_),
    .C(_00646_),
    .Y(_00285_)
  );
  NOR2X1 _06799_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(dbg_0.dbg_rd_rdy ),
    .Y(_00647_)
  );
  NOR2X1 _06800_ (
    .A(_00369_),
    .B(_00647_),
    .Y(dbg_0.dbg_i2c_0.mem_burst_end )
  );
  AND2X1 _06801_ (
    .A(dbg_0.mem_data_0_ ),
    .B(_00377_),
    .Y(_00144_)
  );
  AND2X1 _06802_ (
    .A(dbg_0.mem_data_1_ ),
    .B(_00377_),
    .Y(_00151_)
  );
  AND2X1 _06803_ (
    .A(dbg_0.mem_data_2_ ),
    .B(_00377_),
    .Y(_00152_)
  );
  AND2X1 _06804_ (
    .A(dbg_0.mem_data_3_ ),
    .B(_00377_),
    .Y(_00153_)
  );
  AND2X1 _06805_ (
    .A(dbg_0.mem_data_4_ ),
    .B(_00377_),
    .Y(_00154_)
  );
  AND2X1 _06806_ (
    .A(dbg_0.mem_data_5_ ),
    .B(_00377_),
    .Y(_00155_)
  );
  AND2X1 _06807_ (
    .A(dbg_0.mem_data_6_ ),
    .B(_00377_),
    .Y(_00156_)
  );
  AND2X1 _06808_ (
    .A(dbg_0.mem_data_7_ ),
    .B(_00377_),
    .Y(_00157_)
  );
  NAND2X1 _06809_ (
    .A(dbg_0.mem_data_0_ ),
    .B(_00376_),
    .Y(_00648_)
  );
  OAI21X1 _06810_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00337_),
    .C(_00648_),
    .Y(_00158_)
  );
  NAND2X1 _06811_ (
    .A(dbg_0.mem_data_1_ ),
    .B(_00376_),
    .Y(_00649_)
  );
  OAI21X1 _06812_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00338_),
    .C(_00649_),
    .Y(_00159_)
  );
  NAND2X1 _06813_ (
    .A(dbg_0.mem_data_2_ ),
    .B(_00376_),
    .Y(_00650_)
  );
  OAI21X1 _06814_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00339_),
    .C(_00650_),
    .Y(_00145_)
  );
  NAND2X1 _06815_ (
    .A(dbg_0.mem_data_3_ ),
    .B(_00376_),
    .Y(_00651_)
  );
  OAI21X1 _06816_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00340_),
    .C(_00651_),
    .Y(_00146_)
  );
  NAND2X1 _06817_ (
    .A(dbg_0.mem_data_4_ ),
    .B(_00376_),
    .Y(_00652_)
  );
  OAI21X1 _06818_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00341_),
    .C(_00652_),
    .Y(_00147_)
  );
  NAND2X1 _06819_ (
    .A(dbg_0.mem_data_5_ ),
    .B(_00376_),
    .Y(_00653_)
  );
  OAI21X1 _06820_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00342_),
    .C(_00653_),
    .Y(_00148_)
  );
  NAND2X1 _06821_ (
    .A(dbg_0.mem_data_6_ ),
    .B(_00376_),
    .Y(_00654_)
  );
  OAI21X1 _06822_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00343_),
    .C(_00654_),
    .Y(_00149_)
  );
  NAND2X1 _06823_ (
    .A(dbg_0.mem_data_7_ ),
    .B(_00376_),
    .Y(_00655_)
  );
  OAI21X1 _06824_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00344_),
    .C(_00655_),
    .Y(_00150_)
  );
  AOI21X1 _06825_ (
    .A(_00331_),
    .B(_00577_),
    .C(dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00278_)
  );
  AND2X1 _06826_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(_00385_),
    .Y(_00314_)
  );
  NOR2X1 _06827_ (
    .A(_00328_),
    .B(_00422_),
    .Y(dbg_0.dbg_reg_wr )
  );
  NOR2X1 _06828_ (
    .A(_00392_),
    .B(_00514_),
    .Y(_00656_)
  );
  NOR2X1 _06829_ (
    .A(_00379_),
    .B(_00392_),
    .Y(_00657_)
  );
  OR2X1 _06830_ (
    .A(dbg_0.dbg_addr_5_ ),
    .B(_00379_),
    .Y(_00658_)
  );
  NAND3X1 _06831_ (
    .A(dbg_0.dbg_addr_3_ ),
    .B(dbg_0.dbg_addr_4_ ),
    .C(_00383_),
    .Y(_00659_)
  );
  NOR2X1 _06832_ (
    .A(_00658_),
    .B(_00659_),
    .Y(_00660_)
  );
  AOI22X1 _06833_ (
    .A(dbg_0.mem_data_0_ ),
    .B(_00419_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_0_ ),
    .Y(_00661_)
  );
  INVX1 _06834_ (
    .A(_00661_),
    .Y(_00662_)
  );
  AOI21X1 _06835_ (
    .A(cpu_halt_st),
    .B(_00393_),
    .C(_00662_),
    .Y(_00663_)
  );
  AOI22X1 _06836_ (
    .A(1'h1),
    .B(_00657_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00664_)
  );
  AOI22X1 _06837_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .B(_00515_),
    .C(_00656_),
    .D(1'h1),
    .Y(_00665_)
  );
  NAND3X1 _06838_ (
    .A(_00663_),
    .B(_00664_),
    .C(_00665_),
    .Y(dbg_0.dbg_dout_0_ )
  );
  AOI22X1 _06839_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00384_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00666_)
  );
  AOI22X1 _06840_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .B(_00515_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_1_ ),
    .Y(_00667_)
  );
  AOI22X1 _06841_ (
    .A(1'h0),
    .B(_00656_),
    .C(_00657_),
    .D(1'h1),
    .Y(_00668_)
  );
  INVX1 _06842_ (
    .A(_00668_),
    .Y(_00669_)
  );
  AOI21X1 _06843_ (
    .A(dbg_0.mem_data_1_ ),
    .B(_00419_),
    .C(_00669_),
    .Y(_00670_)
  );
  NAND3X1 _06844_ (
    .A(_00666_),
    .B(_00667_),
    .C(_00670_),
    .Y(dbg_0.dbg_dout_1_ )
  );
  NAND2X1 _06845_ (
    .A(1'h0),
    .B(_00656_),
    .Y(_00671_)
  );
  AOI22X1 _06846_ (
    .A(dbg_0.mem_cnt_2_ ),
    .B(_00581_),
    .C(_00657_),
    .D(1'h0),
    .Y(_00672_)
  );
  AOI22X1 _06847_ (
    .A(dbg_0.dbg_mem_addr_2_ ),
    .B(_00515_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00673_)
  );
  AOI22X1 _06848_ (
    .A(dbg_0.mem_ctl_2_ ),
    .B(_00384_),
    .C(_00393_),
    .D(dbg_0.cpu_stat_2_ ),
    .Y(_00674_)
  );
  NAND2X1 _06849_ (
    .A(_00673_),
    .B(_00674_),
    .Y(_00675_)
  );
  AOI21X1 _06850_ (
    .A(dbg_0.mem_data_2_ ),
    .B(_00419_),
    .C(_00675_),
    .Y(_00676_)
  );
  NAND3X1 _06851_ (
    .A(_00671_),
    .B(_00672_),
    .C(_00676_),
    .Y(dbg_0.dbg_dout_2_ )
  );
  AOI22X1 _06852_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00384_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00677_)
  );
  AOI22X1 _06853_ (
    .A(1'h0),
    .B(_00656_),
    .C(_00657_),
    .D(1'h0),
    .Y(_00678_)
  );
  AOI22X1 _06854_ (
    .A(dbg_0.cpu_stat_3_ ),
    .B(_00393_),
    .C(_00515_),
    .D(dbg_0.dbg_mem_addr_3_ ),
    .Y(_00679_)
  );
  AOI22X1 _06855_ (
    .A(dbg_0.cpu_ctl_3_ ),
    .B(_00413_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_3_ ),
    .Y(_00680_)
  );
  NAND2X1 _06856_ (
    .A(_00679_),
    .B(_00680_),
    .Y(_00681_)
  );
  AOI21X1 _06857_ (
    .A(dbg_0.mem_data_3_ ),
    .B(_00419_),
    .C(_00681_),
    .Y(_00682_)
  );
  NAND3X1 _06858_ (
    .A(_00677_),
    .B(_00678_),
    .C(_00682_),
    .Y(dbg_0.dbg_dout_3_ )
  );
  AOI22X1 _06859_ (
    .A(dbg_0.mem_data_4_ ),
    .B(_00419_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00683_)
  );
  INVX1 _06860_ (
    .A(_00683_),
    .Y(_00684_)
  );
  AOI21X1 _06861_ (
    .A(1'h0),
    .B(_00656_),
    .C(_00684_),
    .Y(_00685_)
  );
  AOI22X1 _06862_ (
    .A(dbg_0.cpu_ctl_4_ ),
    .B(_00413_),
    .C(_00657_),
    .D(1'h0),
    .Y(_00686_)
  );
  AOI22X1 _06863_ (
    .A(dbg_0.dbg_mem_addr_4_ ),
    .B(_00515_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_4_ ),
    .Y(_00687_)
  );
  NAND3X1 _06864_ (
    .A(_00685_),
    .B(_00686_),
    .C(_00687_),
    .Y(dbg_0.dbg_dout_4_ )
  );
  AOI22X1 _06865_ (
    .A(1'h0),
    .B(_00657_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00688_)
  );
  INVX1 _06866_ (
    .A(_00688_),
    .Y(_00689_)
  );
  AOI21X1 _06867_ (
    .A(1'h0),
    .B(_00656_),
    .C(_00689_),
    .Y(_00690_)
  );
  AOI22X1 _06868_ (
    .A(dbg_0.mem_data_5_ ),
    .B(_00419_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_5_ ),
    .Y(_00691_)
  );
  AOI22X1 _06869_ (
    .A(dbg_0.cpu_ctl_5_ ),
    .B(_00413_),
    .C(_00515_),
    .D(dbg_0.dbg_mem_addr_5_ ),
    .Y(_00692_)
  );
  NAND3X1 _06870_ (
    .A(_00690_),
    .B(_00691_),
    .C(_00692_),
    .Y(dbg_0.dbg_dout_5_ )
  );
  AOI22X1 _06871_ (
    .A(dbg_0.mem_data_6_ ),
    .B(_00419_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_6_ ),
    .Y(_00693_)
  );
  INVX1 _06872_ (
    .A(_00693_),
    .Y(_00694_)
  );
  AOI21X1 _06873_ (
    .A(clock_module_0.dbg_cpu_reset ),
    .B(_00413_),
    .C(_00694_),
    .Y(_00695_)
  );
  AOI22X1 _06874_ (
    .A(1'h0),
    .B(_00656_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00696_)
  );
  AOI22X1 _06875_ (
    .A(dbg_0.dbg_mem_addr_6_ ),
    .B(_00515_),
    .C(_00657_),
    .D(1'h0),
    .Y(_00697_)
  );
  NAND3X1 _06876_ (
    .A(_00695_),
    .B(_00696_),
    .C(_00697_),
    .Y(dbg_0.dbg_dout_6_ )
  );
  NAND2X1 _06877_ (
    .A(1'h0),
    .B(_00660_),
    .Y(_00698_)
  );
  AOI22X1 _06878_ (
    .A(dbg_0.dbg_mem_addr_7_ ),
    .B(_00515_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_7_ ),
    .Y(_00699_)
  );
  AOI22X1 _06879_ (
    .A(1'h0),
    .B(_00656_),
    .C(_00657_),
    .D(1'h0),
    .Y(_00700_)
  );
  INVX1 _06880_ (
    .A(_00700_),
    .Y(_00701_)
  );
  AOI21X1 _06881_ (
    .A(dbg_0.mem_data_7_ ),
    .B(_00419_),
    .C(_00701_),
    .Y(_00702_)
  );
  NAND3X1 _06882_ (
    .A(_00698_),
    .B(_00699_),
    .C(_00702_),
    .Y(dbg_0.dbg_dout_7_ )
  );
  NAND2X1 _06883_ (
    .A(1'h1),
    .B(_00656_),
    .Y(_00703_)
  );
  AOI22X1 _06884_ (
    .A(dbg_0.dbg_mem_addr_8_ ),
    .B(_00515_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00704_)
  );
  AOI22X1 _06885_ (
    .A(dbg_0.mem_data_8_ ),
    .B(_00419_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_8_ ),
    .Y(_00705_)
  );
  INVX1 _06886_ (
    .A(_00705_),
    .Y(_00706_)
  );
  AOI21X1 _06887_ (
    .A(1'h0),
    .B(_00657_),
    .C(_00706_),
    .Y(_00707_)
  );
  NAND3X1 _06888_ (
    .A(_00703_),
    .B(_00704_),
    .C(_00707_),
    .Y(dbg_0.dbg_dout_8_ )
  );
  NAND2X1 _06889_ (
    .A(1'h0),
    .B(_00660_),
    .Y(_00708_)
  );
  AOI22X1 _06890_ (
    .A(dbg_0.mem_cnt_9_ ),
    .B(_00581_),
    .C(_00656_),
    .D(1'h0),
    .Y(_00709_)
  );
  AOI22X1 _06891_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .B(_00515_),
    .C(_00657_),
    .D(1'h0),
    .Y(_00710_)
  );
  INVX1 _06892_ (
    .A(_00710_),
    .Y(_00711_)
  );
  AOI21X1 _06893_ (
    .A(dbg_0.mem_data_9_ ),
    .B(_00419_),
    .C(_00711_),
    .Y(_00712_)
  );
  NAND3X1 _06894_ (
    .A(_00708_),
    .B(_00709_),
    .C(_00712_),
    .Y(dbg_0.dbg_dout_9_ )
  );
  NAND2X1 _06895_ (
    .A(1'h0),
    .B(_00660_),
    .Y(_00713_)
  );
  AOI22X1 _06896_ (
    .A(dbg_0.dbg_mem_addr_10_ ),
    .B(_00515_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_10_ ),
    .Y(_00714_)
  );
  AOI22X1 _06897_ (
    .A(1'h0),
    .B(_00656_),
    .C(_00657_),
    .D(1'h0),
    .Y(_00715_)
  );
  INVX1 _06898_ (
    .A(_00715_),
    .Y(_00716_)
  );
  AOI21X1 _06899_ (
    .A(dbg_0.mem_data_10_ ),
    .B(_00419_),
    .C(_00716_),
    .Y(_00717_)
  );
  NAND3X1 _06900_ (
    .A(_00713_),
    .B(_00714_),
    .C(_00717_),
    .Y(dbg_0.dbg_dout_10_ )
  );
  AOI22X1 _06901_ (
    .A(dbg_0.dbg_mem_addr_11_ ),
    .B(_00515_),
    .C(_00656_),
    .D(1'h0),
    .Y(_00718_)
  );
  INVX1 _06902_ (
    .A(_00718_),
    .Y(_00719_)
  );
  AOI21X1 _06903_ (
    .A(1'h0),
    .B(_00657_),
    .C(_00719_),
    .Y(_00720_)
  );
  NAND2X1 _06904_ (
    .A(dbg_0.mem_data_11_ ),
    .B(_00419_),
    .Y(_00721_)
  );
  AOI22X1 _06905_ (
    .A(dbg_0.mem_cnt_11_ ),
    .B(_00581_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00722_)
  );
  NAND3X1 _06906_ (
    .A(_00720_),
    .B(_00721_),
    .C(_00722_),
    .Y(dbg_0.dbg_dout_11_ )
  );
  NAND2X1 _06907_ (
    .A(1'h0),
    .B(_00656_),
    .Y(_00723_)
  );
  AOI22X1 _06908_ (
    .A(dbg_0.dbg_mem_addr_12_ ),
    .B(_00515_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00724_)
  );
  AOI22X1 _06909_ (
    .A(dbg_0.mem_data_12_ ),
    .B(_00419_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_12_ ),
    .Y(_00725_)
  );
  INVX1 _06910_ (
    .A(_00725_),
    .Y(_00726_)
  );
  AOI21X1 _06911_ (
    .A(1'h0),
    .B(_00657_),
    .C(_00726_),
    .Y(_00727_)
  );
  NAND3X1 _06912_ (
    .A(_00723_),
    .B(_00724_),
    .C(_00727_),
    .Y(dbg_0.dbg_dout_12_ )
  );
  NAND2X1 _06913_ (
    .A(1'h0),
    .B(_00660_),
    .Y(_00728_)
  );
  AOI22X1 _06914_ (
    .A(dbg_0.mem_data_13_ ),
    .B(_00419_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_13_ ),
    .Y(_00729_)
  );
  AOI22X1 _06915_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .B(_00515_),
    .C(_00656_),
    .D(1'h0),
    .Y(_00730_)
  );
  INVX1 _06916_ (
    .A(_00730_),
    .Y(_00731_)
  );
  AOI21X1 _06917_ (
    .A(1'h0),
    .B(_00657_),
    .C(_00731_),
    .Y(_00732_)
  );
  NAND3X1 _06918_ (
    .A(_00728_),
    .B(_00729_),
    .C(_00732_),
    .Y(dbg_0.dbg_dout_13_ )
  );
  NAND2X1 _06919_ (
    .A(1'h0),
    .B(_00660_),
    .Y(_00733_)
  );
  AOI22X1 _06920_ (
    .A(dbg_0.dbg_mem_addr_14_ ),
    .B(_00515_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_14_ ),
    .Y(_00734_)
  );
  AOI22X1 _06921_ (
    .A(1'h0),
    .B(_00656_),
    .C(_00657_),
    .D(1'h1),
    .Y(_00735_)
  );
  INVX1 _06922_ (
    .A(_00735_),
    .Y(_00736_)
  );
  AOI21X1 _06923_ (
    .A(dbg_0.mem_data_14_ ),
    .B(_00419_),
    .C(_00736_),
    .Y(_00737_)
  );
  NAND3X1 _06924_ (
    .A(_00733_),
    .B(_00734_),
    .C(_00737_),
    .Y(dbg_0.dbg_dout_14_ )
  );
  NAND2X1 _06925_ (
    .A(1'h1),
    .B(_00656_),
    .Y(_00738_)
  );
  AOI22X1 _06926_ (
    .A(dbg_0.dbg_mem_addr_15_ ),
    .B(_00515_),
    .C(_00660_),
    .D(1'h0),
    .Y(_00739_)
  );
  AOI22X1 _06927_ (
    .A(dbg_0.mem_data_15_ ),
    .B(_00419_),
    .C(_00581_),
    .D(dbg_0.mem_cnt_15_ ),
    .Y(_00740_)
  );
  INVX1 _06928_ (
    .A(_00740_),
    .Y(_00741_)
  );
  AOI21X1 _06929_ (
    .A(1'h0),
    .B(_00657_),
    .C(_00741_),
    .Y(_00742_)
  );
  NAND3X1 _06930_ (
    .A(_00738_),
    .B(_00739_),
    .C(_00742_),
    .Y(dbg_0.dbg_dout_15_ )
  );
  OAI21X1 _06931_ (
    .A(dbg_0.cpu_ctl_4_ ),
    .B(_00355_),
    .C(cpu_halt_st),
    .Y(_00743_)
  );
  INVX1 _06932_ (
    .A(_00743_),
    .Y(_00049_)
  );
  NOR2X1 _06933_ (
    .A(dbg_0.inc_step_1_ ),
    .B(_00511_),
    .Y(cpu_halt_cmd)
  );
  NOR2X1 _06934_ (
    .A(_00328_),
    .B(_00577_),
    .Y(dbg_0.dbg_i2c_0.mem_burst_wr )
  );
  OAI21X1 _06935_ (
    .A(dbg_0.dbg_i2c_0.dbg_wr ),
    .B(dbg_0.dbg_i2c_0.dbg_rd ),
    .C(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00744_)
  );
  OAI21X1 _06936_ (
    .A(dbg_0.mem_ctl_1_ ),
    .B(_00577_),
    .C(_00744_),
    .Y(_00315_)
  );
  AND2X1 _06937_ (
    .A(_00328_),
    .B(dbg_0.dbg_mem_en ),
    .Y(dbg_0.dbg_mem_rd )
  );
  DFFSR _06938_ (
    .CLK(dco_clk),
    .D(_00318_),
    .Q(dbg_0.mem_state_0_ ),
    .R(1'h1),
    .S(_00320_)
  );
  DFFSR _06939_ (
    .CLK(dco_clk),
    .D(_00316_),
    .Q(dbg_0.mem_state_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06940_ (
    .CLK(dco_clk),
    .D(_00319_),
    .Q(dbg_0.mem_state_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06941_ (
    .CLK(dco_clk),
    .D(_00317_),
    .Q(dbg_0.mem_state_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06942_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_mem_rd ),
    .Q(dbg_0.dbg_mem_rd_dly ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06943_ (
    .CLK(dco_clk),
    .D(_00315_),
    .Q(dbg_0.mem_startb ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06944_ (
    .CLK(dco_clk),
    .D(_00278_),
    .Q(dbg_0.dbg_i2c_0.mem_burst ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06945_ (
    .CLK(dco_clk),
    .D(_00260_),
    .Q(dbg_0.halt_flag ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06946_ (
    .CLK(dco_clk),
    .D(dbg_0.istep ),
    .Q(dbg_0.inc_step_0_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06947_ (
    .CLK(dco_clk),
    .D(_00261_),
    .Q(dbg_0.inc_step_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06948_ (
    .CLK(dco_clk),
    .D(_00259_),
    .Q(dbg_0.dbg_rd_rdy ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06949_ (
    .CLK(dco_clk),
    .D(_00279_),
    .Q(dbg_0.mem_cnt_0_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06950_ (
    .CLK(dco_clk),
    .D(_00286_),
    .Q(dbg_0.mem_cnt_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06951_ (
    .CLK(dco_clk),
    .D(_00287_),
    .Q(dbg_0.mem_cnt_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06952_ (
    .CLK(dco_clk),
    .D(_00288_),
    .Q(dbg_0.mem_cnt_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06953_ (
    .CLK(dco_clk),
    .D(_00289_),
    .Q(dbg_0.mem_cnt_4_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06954_ (
    .CLK(dco_clk),
    .D(_00290_),
    .Q(dbg_0.mem_cnt_5_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06955_ (
    .CLK(dco_clk),
    .D(_00291_),
    .Q(dbg_0.mem_cnt_6_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06956_ (
    .CLK(dco_clk),
    .D(_00292_),
    .Q(dbg_0.mem_cnt_7_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06957_ (
    .CLK(dco_clk),
    .D(_00293_),
    .Q(dbg_0.mem_cnt_8_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06958_ (
    .CLK(dco_clk),
    .D(_00294_),
    .Q(dbg_0.mem_cnt_9_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06959_ (
    .CLK(dco_clk),
    .D(_00280_),
    .Q(dbg_0.mem_cnt_10_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06960_ (
    .CLK(dco_clk),
    .D(_00281_),
    .Q(dbg_0.mem_cnt_11_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06961_ (
    .CLK(dco_clk),
    .D(_00282_),
    .Q(dbg_0.mem_cnt_12_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06962_ (
    .CLK(dco_clk),
    .D(_00283_),
    .Q(dbg_0.mem_cnt_13_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06963_ (
    .CLK(dco_clk),
    .D(_00284_),
    .Q(dbg_0.mem_cnt_14_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06964_ (
    .CLK(dco_clk),
    .D(_00285_),
    .Q(dbg_0.mem_cnt_15_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06965_ (
    .CLK(dco_clk),
    .D(_00262_),
    .Q(dbg_0.dbg_mem_addr_0_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06966_ (
    .CLK(dco_clk),
    .D(_00269_),
    .Q(dbg_0.dbg_mem_addr_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06967_ (
    .CLK(dco_clk),
    .D(_00270_),
    .Q(dbg_0.dbg_mem_addr_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06968_ (
    .CLK(dco_clk),
    .D(_00271_),
    .Q(dbg_0.dbg_mem_addr_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06969_ (
    .CLK(dco_clk),
    .D(_00272_),
    .Q(dbg_0.dbg_mem_addr_4_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06970_ (
    .CLK(dco_clk),
    .D(_00273_),
    .Q(dbg_0.dbg_mem_addr_5_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06971_ (
    .CLK(dco_clk),
    .D(_00274_),
    .Q(dbg_0.dbg_mem_addr_6_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06972_ (
    .CLK(dco_clk),
    .D(_00275_),
    .Q(dbg_0.dbg_mem_addr_7_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06973_ (
    .CLK(dco_clk),
    .D(_00276_),
    .Q(dbg_0.dbg_mem_addr_8_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06974_ (
    .CLK(dco_clk),
    .D(_00277_),
    .Q(dbg_0.dbg_mem_addr_9_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06975_ (
    .CLK(dco_clk),
    .D(_00263_),
    .Q(dbg_0.dbg_mem_addr_10_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06976_ (
    .CLK(dco_clk),
    .D(_00264_),
    .Q(dbg_0.dbg_mem_addr_11_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06977_ (
    .CLK(dco_clk),
    .D(_00265_),
    .Q(dbg_0.dbg_mem_addr_12_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06978_ (
    .CLK(dco_clk),
    .D(_00266_),
    .Q(dbg_0.dbg_mem_addr_13_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06979_ (
    .CLK(dco_clk),
    .D(_00267_),
    .Q(dbg_0.dbg_mem_addr_14_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06980_ (
    .CLK(dco_clk),
    .D(_00268_),
    .Q(dbg_0.dbg_mem_addr_15_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06981_ (
    .CLK(dco_clk),
    .D(_00298_),
    .Q(dbg_0.mem_data_0_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06982_ (
    .CLK(dco_clk),
    .D(_00305_),
    .Q(dbg_0.mem_data_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06983_ (
    .CLK(dco_clk),
    .D(_00306_),
    .Q(dbg_0.mem_data_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06984_ (
    .CLK(dco_clk),
    .D(_00307_),
    .Q(dbg_0.mem_data_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06985_ (
    .CLK(dco_clk),
    .D(_00308_),
    .Q(dbg_0.mem_data_4_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06986_ (
    .CLK(dco_clk),
    .D(_00309_),
    .Q(dbg_0.mem_data_5_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06987_ (
    .CLK(dco_clk),
    .D(_00310_),
    .Q(dbg_0.mem_data_6_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06988_ (
    .CLK(dco_clk),
    .D(_00311_),
    .Q(dbg_0.mem_data_7_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06989_ (
    .CLK(dco_clk),
    .D(_00312_),
    .Q(dbg_0.mem_data_8_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06990_ (
    .CLK(dco_clk),
    .D(_00313_),
    .Q(dbg_0.mem_data_9_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06991_ (
    .CLK(dco_clk),
    .D(_00299_),
    .Q(dbg_0.mem_data_10_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06992_ (
    .CLK(dco_clk),
    .D(_00300_),
    .Q(dbg_0.mem_data_11_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06993_ (
    .CLK(dco_clk),
    .D(_00301_),
    .Q(dbg_0.mem_data_12_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06994_ (
    .CLK(dco_clk),
    .D(_00302_),
    .Q(dbg_0.mem_data_13_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06995_ (
    .CLK(dco_clk),
    .D(_00303_),
    .Q(dbg_0.mem_data_14_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06996_ (
    .CLK(dco_clk),
    .D(_00304_),
    .Q(dbg_0.mem_data_15_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06997_ (
    .CLK(dco_clk),
    .D(_00314_),
    .Q(dbg_0.mem_start ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06998_ (
    .CLK(dco_clk),
    .D(_00295_),
    .Q(dbg_0.mem_ctl_1_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _06999_ (
    .CLK(dco_clk),
    .D(_00296_),
    .Q(dbg_0.mem_ctl_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07000_ (
    .CLK(dco_clk),
    .D(_00297_),
    .Q(dbg_0.dbg_i2c_0.mem_bw ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07001_ (
    .CLK(dco_clk),
    .D(_00257_),
    .Q(dbg_0.cpu_stat_2_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07002_ (
    .CLK(dco_clk),
    .D(_00258_),
    .Q(dbg_0.cpu_stat_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07003_ (
    .CLK(dco_clk),
    .D(_00253_),
    .Q(dbg_0.cpu_ctl_3_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07004_ (
    .CLK(dco_clk),
    .D(_00254_),
    .Q(dbg_0.cpu_ctl_4_ ),
    .R(1'h1),
    .S(_00320_)
  );
  DFFSR _07005_ (
    .CLK(dco_clk),
    .D(_00255_),
    .Q(dbg_0.cpu_ctl_5_ ),
    .R(_00320_),
    .S(1'h1)
  );
  DFFSR _07006_ (
    .CLK(dco_clk),
    .D(_00256_),
    .Q(clock_module_0.dbg_cpu_reset ),
    .R(_00320_),
    .S(1'h1)
  );
  INVX1 _07007_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .Y(_00784_)
  );
  INVX1 _07008_ (
    .A(dbg_0.dbg_i2c_0.sda_in_sync_n ),
    .Y(dbg_0.dbg_i2c_0.sda_in_sync )
  );
  INVX1 _07009_ (
    .A(dbg_0.dbg_i2c_0.scl_sync_n ),
    .Y(dbg_0.dbg_i2c_0.scl_sync )
  );
  INVX1 _07010_ (
    .A(dbg_0.dbg_i2c_0.scl_dly ),
    .Y(_00785_)
  );
  INVX1 _07011_ (
    .A(dbg_0.dbg_i2c_0.sda_in_dly ),
    .Y(_00786_)
  );
  INVX1 _07012_ (
    .A(dbg_0.dbg_i2c_0.i2c_active_seq ),
    .Y(_00787_)
  );
  INVX1 _07013_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .Y(_00788_)
  );
  INVX1 _07014_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .Y(_00789_)
  );
  INVX1 _07015_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .Y(_00790_)
  );
  INVX1 _07016_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .Y(_00791_)
  );
  INVX1 _07017_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .Y(_00792_)
  );
  INVX1 _07018_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .Y(_00793_)
  );
  INVX1 _07019_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_3_ ),
    .Y(_00794_)
  );
  INVX1 _07020_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00795_)
  );
  INVX1 _07021_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_5_ ),
    .Y(_00796_)
  );
  INVX1 _07022_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .Y(_00797_)
  );
  INVX1 _07023_ (
    .A(dbg_i2c_addr_2_),
    .Y(_00798_)
  );
  INVX1 _07024_ (
    .A(dbg_i2c_addr_4_),
    .Y(_00799_)
  );
  INVX1 _07025_ (
    .A(dbg_0.dbg_din_8_ ),
    .Y(_00800_)
  );
  INVX1 _07026_ (
    .A(dbg_0.dbg_din_9_ ),
    .Y(_00801_)
  );
  INVX1 _07027_ (
    .A(dbg_0.dbg_din_10_ ),
    .Y(_00802_)
  );
  INVX1 _07028_ (
    .A(dbg_0.dbg_din_11_ ),
    .Y(_00803_)
  );
  INVX1 _07029_ (
    .A(dbg_0.dbg_din_12_ ),
    .Y(_00804_)
  );
  INVX1 _07030_ (
    .A(dbg_0.dbg_din_13_ ),
    .Y(_00805_)
  );
  INVX1 _07031_ (
    .A(dbg_0.dbg_din_14_ ),
    .Y(_00806_)
  );
  INVX1 _07032_ (
    .A(dbg_0.dbg_din_15_ ),
    .Y(_00807_)
  );
  INVX1 _07033_ (
    .A(dbg_0.dbg_dout_0_ ),
    .Y(_00808_)
  );
  INVX1 _07034_ (
    .A(dbg_0.dbg_dout_1_ ),
    .Y(_00809_)
  );
  INVX1 _07035_ (
    .A(dbg_0.dbg_dout_2_ ),
    .Y(_00810_)
  );
  INVX1 _07036_ (
    .A(dbg_0.dbg_dout_3_ ),
    .Y(_00811_)
  );
  INVX1 _07037_ (
    .A(dbg_0.dbg_dout_4_ ),
    .Y(_00812_)
  );
  INVX1 _07038_ (
    .A(dbg_0.dbg_dout_5_ ),
    .Y(_00813_)
  );
  INVX1 _07039_ (
    .A(dbg_0.dbg_dout_6_ ),
    .Y(_00814_)
  );
  INVX1 _07040_ (
    .A(dbg_0.dbg_dout_7_ ),
    .Y(_00815_)
  );
  INVX1 _07041_ (
    .A(dbg_i2c_scl),
    .Y(dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in )
  );
  INVX1 _07042_ (
    .A(dbg_i2c_sda_in),
    .Y(dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in )
  );
  INVX1 _07043_ (
    .A(clock_module_0.dbg_rst ),
    .Y(_00783_)
  );
  OR2X1 _07044_ (
    .A(dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .Y(_00816_)
  );
  AND2X1 _07045_ (
    .A(dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .Y(_00817_)
  );
  OAI21X1 _07046_ (
    .A(dbg_0.dbg_i2c_0.sda_in_sync ),
    .B(_00817_),
    .C(_00816_),
    .Y(_00818_)
  );
  INVX1 _07047_ (
    .A(_00818_),
    .Y(dbg_0.dbg_i2c_0.sda_in )
  );
  OR2X1 _07048_ (
    .A(dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .Y(_00819_)
  );
  AND2X1 _07049_ (
    .A(dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .Y(_00820_)
  );
  OAI21X1 _07050_ (
    .A(dbg_0.dbg_i2c_0.scl_sync ),
    .B(_00820_),
    .C(_00819_),
    .Y(_00821_)
  );
  INVX1 _07051_ (
    .A(_00821_),
    .Y(dbg_0.dbg_i2c_0.scl )
  );
  NOR3X1 _07052_ (
    .A(dbg_0.dbg_i2c_0.sda_in_dly ),
    .B(_00818_),
    .C(_00821_),
    .Y(_00822_)
  );
  NAND3X1 _07053_ (
    .A(_00786_),
    .B(dbg_0.dbg_i2c_0.sda_in ),
    .C(dbg_0.dbg_i2c_0.scl ),
    .Y(_00823_)
  );
  NOR2X1 _07054_ (
    .A(_00787_),
    .B(_00822_),
    .Y(_00824_)
  );
  NOR3X1 _07055_ (
    .A(_00786_),
    .B(dbg_0.dbg_i2c_0.sda_in ),
    .C(_00821_),
    .Y(_00825_)
  );
  NAND3X1 _07056_ (
    .A(dbg_0.dbg_i2c_0.sda_in_dly ),
    .B(_00818_),
    .C(dbg_0.dbg_i2c_0.scl ),
    .Y(_00826_)
  );
  NOR3X1 _07057_ (
    .A(_00787_),
    .B(_00822_),
    .C(_00825_),
    .Y(_00827_)
  );
  NAND3X1 _07058_ (
    .A(dbg_0.dbg_i2c_0.i2c_active_seq ),
    .B(_00823_),
    .C(_00826_),
    .Y(_00828_)
  );
  NAND2X1 _07059_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .B(_00827_),
    .Y(_00829_)
  );
  NOR2X1 _07060_ (
    .A(_00785_),
    .B(dbg_0.dbg_i2c_0.scl ),
    .Y(_00830_)
  );
  NAND2X1 _07061_ (
    .A(dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00821_),
    .Y(_00831_)
  );
  NOR2X1 _07062_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .Y(_00832_)
  );
  NAND2X1 _07063_ (
    .A(_00793_),
    .B(_00832_),
    .Y(_00833_)
  );
  NAND2X1 _07064_ (
    .A(_00790_),
    .B(_00791_),
    .Y(_00834_)
  );
  NOR2X1 _07065_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .Y(_00835_)
  );
  NAND3X1 _07066_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(_00789_),
    .C(_00835_),
    .Y(_00836_)
  );
  NOR3X1 _07067_ (
    .A(_00833_),
    .B(_00834_),
    .C(_00836_),
    .Y(_00837_)
  );
  NAND2X1 _07068_ (
    .A(_00830_),
    .B(_00837_),
    .Y(_00838_)
  );
  NOR2X1 _07069_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .B(dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .Y(_00839_)
  );
  NOR2X1 _07070_ (
    .A(_00838_),
    .B(_00839_),
    .Y(_00840_)
  );
  NAND2X1 _07071_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(dbg_0.dbg_i2c_0.i2c_state_3_ ),
    .Y(_00841_)
  );
  NAND2X1 _07072_ (
    .A(_00784_),
    .B(_00841_),
    .Y(_00842_)
  );
  OAI21X1 _07073_ (
    .A(_00784_),
    .B(dbg_0.dbg_i2c_0.sda_in ),
    .C(_00841_),
    .Y(_00843_)
  );
  NAND3X1 _07074_ (
    .A(_00824_),
    .B(_00830_),
    .C(_00843_),
    .Y(_00844_)
  );
  OAI21X1 _07075_ (
    .A(_00829_),
    .B(_00840_),
    .C(_00844_),
    .Y(_00778_)
  );
  OAI21X1 _07076_ (
    .A(_00838_),
    .B(_00839_),
    .C(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .Y(_00845_)
  );
  NAND2X1 _07077_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_4_ ),
    .B(_00840_),
    .Y(_00846_)
  );
  NAND2X1 _07078_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(dbg_0.dbg_i2c_0.mem_burst ),
    .Y(_00847_)
  );
  NAND2X1 _07079_ (
    .A(_00795_),
    .B(dbg_0.dbg_i2c_0.dbg_bw ),
    .Y(_00848_)
  );
  AND2X1 _07080_ (
    .A(_00847_),
    .B(_00848_),
    .Y(_00849_)
  );
  INVX1 _07081_ (
    .A(_00849_),
    .Y(_00850_)
  );
  OAI21X1 _07082_ (
    .A(_00846_),
    .B(_00850_),
    .C(_00845_),
    .Y(_00773_)
  );
  NOR3X1 _07083_ (
    .A(_00785_),
    .B(_00788_),
    .C(dbg_0.dbg_i2c_0.scl ),
    .Y(_00851_)
  );
  AND2X1 _07084_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B(_00851_),
    .Y(_00852_)
  );
  NAND2X1 _07085_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B(_00851_),
    .Y(_00853_)
  );
  NAND2X1 _07086_ (
    .A(_00827_),
    .B(_00852_),
    .Y(_00854_)
  );
  OAI21X1 _07087_ (
    .A(_00785_),
    .B(dbg_0.dbg_i2c_0.scl ),
    .C(_00827_),
    .Y(_00855_)
  );
  OAI21X1 _07088_ (
    .A(_00796_),
    .B(_00855_),
    .C(_00854_),
    .Y(_00782_)
  );
  NAND2X1 _07089_ (
    .A(_00796_),
    .B(_00797_),
    .Y(_00856_)
  );
  XOR2X1 _07090_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(dbg_i2c_addr_1_),
    .Y(_00857_)
  );
  XNOR2X1 _07091_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .B(dbg_i2c_addr_0_),
    .Y(_00858_)
  );
  XNOR2X1 _07092_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(dbg_i2c_addr_6_),
    .Y(_00859_)
  );
  XNOR2X1 _07093_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(dbg_i2c_addr_3_),
    .Y(_00860_)
  );
  AOI22X1 _07094_ (
    .A(_00790_),
    .B(dbg_i2c_addr_2_),
    .C(dbg_i2c_addr_4_),
    .D(_00792_),
    .Y(_00861_)
  );
  XOR2X1 _07095_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(dbg_i2c_addr_5_),
    .Y(_00862_)
  );
  AOI22X1 _07096_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(_00798_),
    .C(_00799_),
    .D(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .Y(_00863_)
  );
  NOR2X1 _07097_ (
    .A(_00857_),
    .B(_00862_),
    .Y(_00864_)
  );
  NAND3X1 _07098_ (
    .A(_00859_),
    .B(_00863_),
    .C(_00864_),
    .Y(_00865_)
  );
  NAND3X1 _07099_ (
    .A(_00858_),
    .B(_00860_),
    .C(_00861_),
    .Y(_00866_)
  );
  NOR2X1 _07100_ (
    .A(_00865_),
    .B(_00866_),
    .Y(_00867_)
  );
  AOI21X1 _07101_ (
    .A(_00851_),
    .B(_00867_),
    .C(_00797_),
    .Y(_00868_)
  );
  NAND2X1 _07102_ (
    .A(dbg_0.dbg_i2c_0.sda_in ),
    .B(_00830_),
    .Y(_00869_)
  );
  NOR2X1 _07103_ (
    .A(_00828_),
    .B(_00868_),
    .Y(_00870_)
  );
  OAI21X1 _07104_ (
    .A(_00784_),
    .B(_00869_),
    .C(_00870_),
    .Y(_00777_)
  );
  NOR2X1 _07105_ (
    .A(dbg_0.dbg_i2c_0.mem_burst_rd ),
    .B(dbg_0.dbg_i2c_0.mem_burst_wr ),
    .Y(_00871_)
  );
  AND2X1 _07106_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00852_),
    .Y(_00872_)
  );
  NAND2X1 _07107_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00852_),
    .Y(_00873_)
  );
  NOR2X1 _07108_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(_00873_),
    .Y(_00874_)
  );
  NAND2X1 _07109_ (
    .A(_00871_),
    .B(_00874_),
    .Y(_00875_)
  );
  NAND2X1 _07110_ (
    .A(_00840_),
    .B(_00847_),
    .Y(_00876_)
  );
  NAND2X1 _07111_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00840_),
    .Y(_00877_)
  );
  NAND3X1 _07112_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .C(_00840_),
    .Y(_00878_)
  );
  NAND2X1 _07113_ (
    .A(dbg_0.dbg_i2c_0.mem_burst_rd ),
    .B(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .Y(_00879_)
  );
  OAI21X1 _07114_ (
    .A(dbg_0.dbg_i2c_0.mem_burst_wr ),
    .B(_00879_),
    .C(_00878_),
    .Y(_00880_)
  );
  AOI21X1 _07115_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_4_ ),
    .B(_00876_),
    .C(_00880_),
    .Y(_00881_)
  );
  NAND2X1 _07116_ (
    .A(_00875_),
    .B(_00881_),
    .Y(_00776_)
  );
  NAND3X1 _07117_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .B(_00827_),
    .C(_00831_),
    .Y(_00882_)
  );
  OAI21X1 _07118_ (
    .A(_00829_),
    .B(_00838_),
    .C(_00882_),
    .Y(_00781_)
  );
  NOR2X1 _07119_ (
    .A(_00795_),
    .B(dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00883_)
  );
  NAND2X1 _07120_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .B(_00852_),
    .Y(_00884_)
  );
  INVX1 _07121_ (
    .A(_00884_),
    .Y(_00885_)
  );
  AOI21X1 _07122_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_i2c_0.dbg_state_3_ ),
    .C(_00885_),
    .Y(_00886_)
  );
  NAND2X1 _07123_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_3_ ),
    .B(_00852_),
    .Y(_00887_)
  );
  AOI21X1 _07124_ (
    .A(_00846_),
    .B(_00887_),
    .C(_00848_),
    .Y(_00888_)
  );
  NAND3X1 _07125_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .B(_00853_),
    .C(_00871_),
    .Y(_00889_)
  );
  OAI21X1 _07126_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(_00877_),
    .C(_00889_),
    .Y(_00890_)
  );
  NOR2X1 _07127_ (
    .A(_00888_),
    .B(_00890_),
    .Y(_00891_)
  );
  OAI21X1 _07128_ (
    .A(_00883_),
    .B(_00886_),
    .C(_00891_),
    .Y(_00772_)
  );
  NAND2X1 _07129_ (
    .A(_00847_),
    .B(_00852_),
    .Y(_00892_)
  );
  AND2X1 _07130_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00893_)
  );
  NAND2X1 _07131_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_i2c_0.mem_burst_end ),
    .Y(_00894_)
  );
  NAND2X1 _07132_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(_00871_),
    .Y(_00895_)
  );
  NOR2X1 _07133_ (
    .A(_00853_),
    .B(_00895_),
    .Y(_00896_)
  );
  OAI21X1 _07134_ (
    .A(dbg_0.dbg_i2c_0.mem_burst_wr ),
    .B(_00896_),
    .C(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .Y(_00897_)
  );
  AOI22X1 _07135_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(_00885_),
    .C(_00892_),
    .D(dbg_0.dbg_i2c_0.dbg_state_3_ ),
    .Y(_00898_)
  );
  OAI21X1 _07136_ (
    .A(_00893_),
    .B(_00898_),
    .C(_00897_),
    .Y(_00775_)
  );
  NAND3X1 _07137_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_3_ ),
    .B(_00849_),
    .C(_00894_),
    .Y(_00899_)
  );
  NAND2X1 _07138_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .B(_00853_),
    .Y(_00900_)
  );
  OAI21X1 _07139_ (
    .A(_00853_),
    .B(_00899_),
    .C(_00900_),
    .Y(_00774_)
  );
  AND2X1 _07140_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .B(_00851_),
    .Y(_00901_)
  );
  NAND2X1 _07141_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .B(_00851_),
    .Y(_00902_)
  );
  NAND3X1 _07142_ (
    .A(_00827_),
    .B(_00867_),
    .C(_00901_),
    .Y(_00903_)
  );
  OAI21X1 _07143_ (
    .A(_00794_),
    .B(_00855_),
    .C(_00903_),
    .Y(_00780_)
  );
  OAI21X1 _07144_ (
    .A(_00788_),
    .B(_00831_),
    .C(dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .Y(_00904_)
  );
  OAI21X1 _07145_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00794_),
    .C(_00796_),
    .Y(_00905_)
  );
  NAND2X1 _07146_ (
    .A(_00830_),
    .B(_00905_),
    .Y(_00906_)
  );
  AOI21X1 _07147_ (
    .A(_00904_),
    .B(_00906_),
    .C(_00828_),
    .Y(_00779_)
  );
  NAND2X1 _07148_ (
    .A(_00795_),
    .B(dbg_0.dbg_addr_0_ ),
    .Y(_00907_)
  );
  NAND2X1 _07149_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00872_),
    .Y(_00908_)
  );
  OAI21X1 _07150_ (
    .A(_00872_),
    .B(_00907_),
    .C(_00908_),
    .Y(_00745_)
  );
  OAI21X1 _07151_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_addr_1_ ),
    .C(_00873_),
    .Y(_00909_)
  );
  OAI21X1 _07152_ (
    .A(_00789_),
    .B(_00873_),
    .C(_00909_),
    .Y(_00746_)
  );
  OAI21X1 _07153_ (
    .A(dbg_0.dbg_i2c_0.mem_burst ),
    .B(dbg_0.dbg_addr_2_ ),
    .C(_00873_),
    .Y(_00910_)
  );
  OAI21X1 _07154_ (
    .A(_00791_),
    .B(_00873_),
    .C(_00910_),
    .Y(_00747_)
  );
  AOI21X1 _07155_ (
    .A(_00795_),
    .B(dbg_0.dbg_addr_3_ ),
    .C(_00872_),
    .Y(_00911_)
  );
  AOI21X1 _07156_ (
    .A(_00790_),
    .B(_00872_),
    .C(_00911_),
    .Y(_00748_)
  );
  NAND2X1 _07157_ (
    .A(_00795_),
    .B(dbg_0.dbg_addr_4_ ),
    .Y(_00912_)
  );
  NAND2X1 _07158_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(_00872_),
    .Y(_00913_)
  );
  OAI21X1 _07159_ (
    .A(_00872_),
    .B(_00912_),
    .C(_00913_),
    .Y(_00749_)
  );
  AOI21X1 _07160_ (
    .A(_00795_),
    .B(dbg_0.dbg_addr_5_ ),
    .C(_00872_),
    .Y(_00914_)
  );
  AOI21X1 _07161_ (
    .A(_00792_),
    .B(_00872_),
    .C(_00914_),
    .Y(_00750_)
  );
  NAND2X1 _07162_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(_00872_),
    .Y(_00915_)
  );
  OAI21X1 _07163_ (
    .A(_00849_),
    .B(_00872_),
    .C(_00915_),
    .Y(_00751_)
  );
  OAI21X1 _07164_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00884_),
    .C(_00887_),
    .Y(_00916_)
  );
  AOI21X1 _07165_ (
    .A(_00800_),
    .B(_00884_),
    .C(_00916_),
    .Y(_00752_)
  );
  OAI21X1 _07166_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .B(_00884_),
    .C(_00887_),
    .Y(_00917_)
  );
  AOI21X1 _07167_ (
    .A(_00801_),
    .B(_00884_),
    .C(_00917_),
    .Y(_00753_)
  );
  OAI21X1 _07168_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(_00884_),
    .C(_00887_),
    .Y(_00918_)
  );
  AOI21X1 _07169_ (
    .A(_00802_),
    .B(_00884_),
    .C(_00918_),
    .Y(_00754_)
  );
  OAI21X1 _07170_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(_00884_),
    .C(_00887_),
    .Y(_00919_)
  );
  AOI21X1 _07171_ (
    .A(_00803_),
    .B(_00884_),
    .C(_00919_),
    .Y(_00755_)
  );
  OAI21X1 _07172_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(_00884_),
    .C(_00887_),
    .Y(_00920_)
  );
  AOI21X1 _07173_ (
    .A(_00804_),
    .B(_00884_),
    .C(_00920_),
    .Y(_00756_)
  );
  OAI21X1 _07174_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(_00884_),
    .C(_00887_),
    .Y(_00921_)
  );
  AOI21X1 _07175_ (
    .A(_00805_),
    .B(_00884_),
    .C(_00921_),
    .Y(_00757_)
  );
  OAI21X1 _07176_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(_00884_),
    .C(_00887_),
    .Y(_00922_)
  );
  AOI21X1 _07177_ (
    .A(_00806_),
    .B(_00884_),
    .C(_00922_),
    .Y(_00758_)
  );
  OAI21X1 _07178_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(_00884_),
    .C(_00887_),
    .Y(_00923_)
  );
  AOI21X1 _07179_ (
    .A(_00807_),
    .B(_00884_),
    .C(_00923_),
    .Y(_00759_)
  );
  MUX2X1 _07180_ (
    .A(dbg_0.dbg_din_0_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .S(_00887_),
    .Y(_00924_)
  );
  INVX1 _07181_ (
    .A(_00924_),
    .Y(_00760_)
  );
  MUX2X1 _07182_ (
    .A(dbg_0.dbg_din_1_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .S(_00887_),
    .Y(_00925_)
  );
  INVX1 _07183_ (
    .A(_00925_),
    .Y(_00761_)
  );
  MUX2X1 _07184_ (
    .A(dbg_0.dbg_din_2_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .S(_00887_),
    .Y(_00926_)
  );
  INVX1 _07185_ (
    .A(_00926_),
    .Y(_00762_)
  );
  MUX2X1 _07186_ (
    .A(dbg_0.dbg_din_3_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .S(_00887_),
    .Y(_00927_)
  );
  INVX1 _07187_ (
    .A(_00927_),
    .Y(_00763_)
  );
  MUX2X1 _07188_ (
    .A(dbg_0.dbg_din_4_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .S(_00887_),
    .Y(_00928_)
  );
  INVX1 _07189_ (
    .A(_00928_),
    .Y(_00764_)
  );
  MUX2X1 _07190_ (
    .A(dbg_0.dbg_din_5_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .S(_00887_),
    .Y(_00929_)
  );
  INVX1 _07191_ (
    .A(_00929_),
    .Y(_00765_)
  );
  MUX2X1 _07192_ (
    .A(dbg_0.dbg_din_6_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .S(_00887_),
    .Y(_00930_)
  );
  INVX1 _07193_ (
    .A(_00930_),
    .Y(_00766_)
  );
  MUX2X1 _07194_ (
    .A(dbg_0.dbg_din_7_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .S(_00887_),
    .Y(_00931_)
  );
  INVX1 _07195_ (
    .A(_00931_),
    .Y(_00767_)
  );
  OAI21X1 _07196_ (
    .A(_00785_),
    .B(dbg_0.dbg_i2c_0.scl ),
    .C(_00050_),
    .Y(_00932_)
  );
  NAND3X1 _07197_ (
    .A(_00829_),
    .B(_00844_),
    .C(_00882_),
    .Y(_00933_)
  );
  NOR2X1 _07198_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_3_ ),
    .B(dbg_0.dbg_i2c_0.i2c_state_5_ ),
    .Y(_00934_)
  );
  AOI21X1 _07199_ (
    .A(_00784_),
    .B(_00934_),
    .C(_00855_),
    .Y(_00935_)
  );
  OAI21X1 _07200_ (
    .A(_00829_),
    .B(_00838_),
    .C(_00903_),
    .Y(_00936_)
  );
  NOR2X1 _07201_ (
    .A(_00935_),
    .B(_00936_),
    .Y(_00937_)
  );
  AOI21X1 _07202_ (
    .A(_00854_),
    .B(_00937_),
    .C(_00933_),
    .Y(_00938_)
  );
  NOR2X1 _07203_ (
    .A(_00831_),
    .B(_00837_),
    .Y(_00939_)
  );
  OAI21X1 _07204_ (
    .A(_00828_),
    .B(_00853_),
    .C(_00939_),
    .Y(_00940_)
  );
  NOR2X1 _07205_ (
    .A(_00779_),
    .B(_00940_),
    .Y(_00941_)
  );
  OAI21X1 _07206_ (
    .A(_00778_),
    .B(_00781_),
    .C(_00941_),
    .Y(_00942_)
  );
  OAI21X1 _07207_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(_00942_),
    .C(_00830_),
    .Y(_00943_)
  );
  OAI21X1 _07208_ (
    .A(_00938_),
    .B(_00943_),
    .C(_00932_),
    .Y(_00768_)
  );
  NOR2X1 _07209_ (
    .A(dbg_0.dbg_i2c_0.scl_dly ),
    .B(_00821_),
    .Y(dbg_0.dbg_i2c_0.scl_re )
  );
  OAI21X1 _07210_ (
    .A(dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .B(_00856_),
    .C(dbg_0.dbg_i2c_0.scl_re_dly_1_ ),
    .Y(_00944_)
  );
  INVX1 _07211_ (
    .A(_00944_),
    .Y(_00945_)
  );
  AOI21X1 _07212_ (
    .A(_00933_),
    .B(_00941_),
    .C(_00945_),
    .Y(_00946_)
  );
  NAND2X1 _07213_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .B(_00946_),
    .Y(_00947_)
  );
  AND2X1 _07214_ (
    .A(_00827_),
    .B(_00906_),
    .Y(_00948_)
  );
  NAND2X1 _07215_ (
    .A(_00842_),
    .B(dbg_0.dbg_i2c_0.scl_re ),
    .Y(_00949_)
  );
  OAI21X1 _07216_ (
    .A(_00818_),
    .B(_00944_),
    .C(_00948_),
    .Y(_00950_)
  );
  INVX1 _07217_ (
    .A(_00950_),
    .Y(_00951_)
  );
  NAND3X1 _07218_ (
    .A(_00947_),
    .B(_00949_),
    .C(_00951_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_0_ )
  );
  MUX2X1 _07219_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .S(_00946_),
    .Y(_00952_)
  );
  NAND2X1 _07220_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_8_ ),
    .Y(_00953_)
  );
  OAI21X1 _07221_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00808_),
    .C(_00953_),
    .Y(_00954_)
  );
  OAI21X1 _07222_ (
    .A(_00949_),
    .B(_00954_),
    .C(_00948_),
    .Y(_00955_)
  );
  AOI21X1 _07223_ (
    .A(_00949_),
    .B(_00952_),
    .C(_00955_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_1_ )
  );
  MUX2X1 _07224_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .S(_00946_),
    .Y(_00956_)
  );
  NAND2X1 _07225_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_9_ ),
    .Y(_00957_)
  );
  OAI21X1 _07226_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00809_),
    .C(_00957_),
    .Y(_00958_)
  );
  OAI21X1 _07227_ (
    .A(_00949_),
    .B(_00958_),
    .C(_00948_),
    .Y(_00959_)
  );
  AOI21X1 _07228_ (
    .A(_00949_),
    .B(_00956_),
    .C(_00959_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_2_ )
  );
  MUX2X1 _07229_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .S(_00946_),
    .Y(_00960_)
  );
  NAND2X1 _07230_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_10_ ),
    .Y(_00961_)
  );
  OAI21X1 _07231_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00810_),
    .C(_00961_),
    .Y(_00962_)
  );
  OAI21X1 _07232_ (
    .A(_00949_),
    .B(_00962_),
    .C(_00948_),
    .Y(_00963_)
  );
  AOI21X1 _07233_ (
    .A(_00949_),
    .B(_00960_),
    .C(_00963_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_3_ )
  );
  MUX2X1 _07234_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .S(_00946_),
    .Y(_00964_)
  );
  NAND2X1 _07235_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_11_ ),
    .Y(_00965_)
  );
  OAI21X1 _07236_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00811_),
    .C(_00965_),
    .Y(_00966_)
  );
  OAI21X1 _07237_ (
    .A(_00949_),
    .B(_00966_),
    .C(_00948_),
    .Y(_00967_)
  );
  AOI21X1 _07238_ (
    .A(_00949_),
    .B(_00964_),
    .C(_00967_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_4_ )
  );
  MUX2X1 _07239_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .S(_00946_),
    .Y(_00968_)
  );
  NAND2X1 _07240_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_12_ ),
    .Y(_00969_)
  );
  OAI21X1 _07241_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00812_),
    .C(_00969_),
    .Y(_00970_)
  );
  OAI21X1 _07242_ (
    .A(_00949_),
    .B(_00970_),
    .C(_00948_),
    .Y(_00971_)
  );
  AOI21X1 _07243_ (
    .A(_00949_),
    .B(_00968_),
    .C(_00971_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_5_ )
  );
  MUX2X1 _07244_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .S(_00946_),
    .Y(_00972_)
  );
  NAND2X1 _07245_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_13_ ),
    .Y(_00973_)
  );
  OAI21X1 _07246_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00813_),
    .C(_00973_),
    .Y(_00974_)
  );
  OAI21X1 _07247_ (
    .A(_00949_),
    .B(_00974_),
    .C(_00948_),
    .Y(_00975_)
  );
  AOI21X1 _07248_ (
    .A(_00949_),
    .B(_00972_),
    .C(_00975_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_6_ )
  );
  MUX2X1 _07249_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .S(_00946_),
    .Y(_00976_)
  );
  NAND2X1 _07250_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_14_ ),
    .Y(_00977_)
  );
  OAI21X1 _07251_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00814_),
    .C(_00977_),
    .Y(_00978_)
  );
  OAI21X1 _07252_ (
    .A(_00949_),
    .B(_00978_),
    .C(_00948_),
    .Y(_00979_)
  );
  AOI21X1 _07253_ (
    .A(_00949_),
    .B(_00976_),
    .C(_00979_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_7_ )
  );
  MUX2X1 _07254_ (
    .A(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .B(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .S(_00946_),
    .Y(_00980_)
  );
  NAND2X1 _07255_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(dbg_0.dbg_dout_15_ ),
    .Y(_00981_)
  );
  OAI21X1 _07256_ (
    .A(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .B(_00815_),
    .C(_00981_),
    .Y(_00982_)
  );
  OAI21X1 _07257_ (
    .A(_00949_),
    .B(_00982_),
    .C(_00948_),
    .Y(_00983_)
  );
  AOI21X1 _07258_ (
    .A(_00949_),
    .B(_00980_),
    .C(_00983_),
    .Y(dbg_0.dbg_i2c_0.shift_buf_nxt_8_ )
  );
  NAND2X1 _07259_ (
    .A(_00849_),
    .B(_00885_),
    .Y(_00984_)
  );
  OAI21X1 _07260_ (
    .A(_00849_),
    .B(_00887_),
    .C(_00984_),
    .Y(_00770_)
  );
  NOR2X1 _07261_ (
    .A(_00846_),
    .B(_00847_),
    .Y(_00985_)
  );
  AOI21X1 _07262_ (
    .A(_00795_),
    .B(_00874_),
    .C(_00985_),
    .Y(_00986_)
  );
  OAI21X1 _07263_ (
    .A(dbg_0.dbg_i2c_0.mem_bw ),
    .B(_00878_),
    .C(_00986_),
    .Y(_00769_)
  );
  OAI21X1 _07264_ (
    .A(_00867_),
    .B(_00902_),
    .C(_00824_),
    .Y(_00987_)
  );
  NAND2X1 _07265_ (
    .A(_00826_),
    .B(_00987_),
    .Y(_00771_)
  );
  DFFSR _07266_ (
    .CLK(dco_clk),
    .D(_00772_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_0_ ),
    .R(1'h1),
    .S(_00783_)
  );
  DFFSR _07267_ (
    .CLK(dco_clk),
    .D(_00773_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_1_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07268_ (
    .CLK(dco_clk),
    .D(_00774_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_2_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07269_ (
    .CLK(dco_clk),
    .D(_00775_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_3_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07270_ (
    .CLK(dco_clk),
    .D(_00776_),
    .Q(dbg_0.dbg_i2c_0.dbg_state_4_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07271_ (
    .CLK(dco_clk),
    .D(_00777_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_0_ ),
    .R(1'h1),
    .S(_00783_)
  );
  DFFSR _07272_ (
    .CLK(dco_clk),
    .D(_00778_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_1_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07273_ (
    .CLK(dco_clk),
    .D(_00779_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_2_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07274_ (
    .CLK(dco_clk),
    .D(_00780_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_3_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07275_ (
    .CLK(dco_clk),
    .D(_00781_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_4_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07276_ (
    .CLK(dco_clk),
    .D(_00782_),
    .Q(dbg_0.dbg_i2c_0.i2c_state_5_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07277_ (
    .CLK(dco_clk),
    .D(_00769_),
    .Q(dbg_0.dbg_i2c_0.dbg_rd ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07278_ (
    .CLK(dco_clk),
    .D(_00770_),
    .Q(dbg_0.dbg_i2c_0.dbg_wr ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07279_ (
    .CLK(dco_clk),
    .D(_00752_),
    .Q(dbg_0.dbg_din_8_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07280_ (
    .CLK(dco_clk),
    .D(_00753_),
    .Q(dbg_0.dbg_din_9_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07281_ (
    .CLK(dco_clk),
    .D(_00754_),
    .Q(dbg_0.dbg_din_10_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07282_ (
    .CLK(dco_clk),
    .D(_00755_),
    .Q(dbg_0.dbg_din_11_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07283_ (
    .CLK(dco_clk),
    .D(_00756_),
    .Q(dbg_0.dbg_din_12_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07284_ (
    .CLK(dco_clk),
    .D(_00757_),
    .Q(dbg_0.dbg_din_13_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07285_ (
    .CLK(dco_clk),
    .D(_00758_),
    .Q(dbg_0.dbg_din_14_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07286_ (
    .CLK(dco_clk),
    .D(_00759_),
    .Q(dbg_0.dbg_din_15_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07287_ (
    .CLK(dco_clk),
    .D(_00760_),
    .Q(dbg_0.dbg_din_0_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07288_ (
    .CLK(dco_clk),
    .D(_00761_),
    .Q(dbg_0.dbg_din_1_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07289_ (
    .CLK(dco_clk),
    .D(_00762_),
    .Q(dbg_0.dbg_din_2_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07290_ (
    .CLK(dco_clk),
    .D(_00763_),
    .Q(dbg_0.dbg_din_3_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07291_ (
    .CLK(dco_clk),
    .D(_00764_),
    .Q(dbg_0.dbg_din_4_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07292_ (
    .CLK(dco_clk),
    .D(_00765_),
    .Q(dbg_0.dbg_din_5_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07293_ (
    .CLK(dco_clk),
    .D(_00766_),
    .Q(dbg_0.dbg_din_6_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07294_ (
    .CLK(dco_clk),
    .D(_00767_),
    .Q(dbg_0.dbg_din_7_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07295_ (
    .CLK(dco_clk),
    .D(_00745_),
    .Q(dbg_0.dbg_addr_0_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07296_ (
    .CLK(dco_clk),
    .D(_00746_),
    .Q(dbg_0.dbg_addr_1_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07297_ (
    .CLK(dco_clk),
    .D(_00747_),
    .Q(dbg_0.dbg_addr_2_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07298_ (
    .CLK(dco_clk),
    .D(_00748_),
    .Q(dbg_0.dbg_addr_3_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07299_ (
    .CLK(dco_clk),
    .D(_00749_),
    .Q(dbg_0.dbg_addr_4_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07300_ (
    .CLK(dco_clk),
    .D(_00750_),
    .Q(dbg_0.dbg_addr_5_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07301_ (
    .CLK(dco_clk),
    .D(_00751_),
    .Q(dbg_0.dbg_i2c_0.dbg_bw ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07302_ (
    .CLK(dco_clk),
    .D(_00768_),
    .Q(_00050_),
    .R(1'h1),
    .S(_00783_)
  );
  DFFSR _07303_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_0_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_0_ ),
    .R(1'h1),
    .S(_00783_)
  );
  DFFSR _07304_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_1_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_1_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07305_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_2_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_2_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07306_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_3_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_3_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07307_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_4_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_4_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07308_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_5_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_5_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07309_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_6_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_6_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07310_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_7_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_7_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07311_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.shift_buf_nxt_8_ ),
    .Q(dbg_0.dbg_i2c_0.shift_buf_8_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07312_ (
    .CLK(dco_clk),
    .D(_00771_),
    .Q(dbg_0.dbg_i2c_0.i2c_active_seq ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07313_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl_re ),
    .Q(dbg_0.dbg_i2c_0.scl_re_dly_0_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07314_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl_re_dly_0_ ),
    .Q(dbg_0.dbg_i2c_0.scl_re_dly_1_ ),
    .R(_00783_),
    .S(1'h1)
  );
  DFFSR _07315_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl ),
    .Q(dbg_0.dbg_i2c_0.scl_dly ),
    .R(1'h1),
    .S(_00783_)
  );
  DFFSR _07316_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sda_in ),
    .Q(dbg_0.dbg_i2c_0.sda_in_dly ),
    .R(1'h1),
    .S(_00783_)
  );
  DFFSR _07317_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sda_in_sync ),
    .Q(dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .R(1'h1),
    .S(_00783_)
  );
  DFFSR _07318_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sda_in_buf_0_ ),
    .Q(dbg_0.dbg_i2c_0.sda_in_buf_1_ ),
    .R(1'h1),
    .S(_00783_)
  );
  DFFSR _07319_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl_sync ),
    .Q(dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .R(1'h1),
    .S(_00783_)
  );
  DFFSR _07320_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.scl_buf_0_ ),
    .Q(dbg_0.dbg_i2c_0.scl_buf_1_ ),
    .R(1'h1),
    .S(_00783_)
  );
  INVX1 _07321_ (
    .A(clock_module_0.dbg_rst ),
    .Y(_00988_)
  );
  DFFSR _07322_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_in ),
    .Q(dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ),
    .R(_00988_),
    .S(1'h1)
  );
  DFFSR _07323_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sync_cell_i2c_scl.data_sync_0_ ),
    .Q(dbg_0.dbg_i2c_0.scl_sync_n ),
    .R(_00988_),
    .S(1'h1)
  );
  INVX1 _07324_ (
    .A(clock_module_0.dbg_rst ),
    .Y(_00989_)
  );
  DFFSR _07325_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_in ),
    .Q(dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ),
    .R(_00989_),
    .S(1'h1)
  );
  DFFSR _07326_ (
    .CLK(dco_clk),
    .D(dbg_0.dbg_i2c_0.sync_cell_i2c_sda.data_sync_0_ ),
    .Q(dbg_0.dbg_i2c_0.sda_in_sync_n ),
    .R(_00989_),
    .S(1'h1)
  );
  INVX1 _07327_ (
    .A(e_state_0_),
    .Y(_01026_)
  );
  INVX1 _07328_ (
    .A(e_state_2_),
    .Y(_01027_)
  );
  INVX1 _07329_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .Y(_01028_)
  );
  INVX1 _07330_ (
    .A(execution_unit_0.mdb_out_nxt_8_ ),
    .Y(_01029_)
  );
  INVX1 _07331_ (
    .A(execution_unit_0.mdb_out_nxt_9_ ),
    .Y(_01030_)
  );
  INVX1 _07332_ (
    .A(execution_unit_0.mdb_out_nxt_10_ ),
    .Y(_01031_)
  );
  INVX1 _07333_ (
    .A(execution_unit_0.mdb_out_nxt_11_ ),
    .Y(_01032_)
  );
  INVX1 _07334_ (
    .A(execution_unit_0.mdb_out_nxt_12_ ),
    .Y(_01033_)
  );
  INVX1 _07335_ (
    .A(execution_unit_0.mdb_out_nxt_13_ ),
    .Y(_01034_)
  );
  INVX1 _07336_ (
    .A(execution_unit_0.mdb_out_nxt_14_ ),
    .Y(_01035_)
  );
  INVX1 _07337_ (
    .A(execution_unit_0.mdb_out_nxt_15_ ),
    .Y(_01036_)
  );
  INVX1 _07338_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_01037_)
  );
  INVX1 _07339_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_alu ),
    .Y(_01038_)
  );
  INVX1 _07340_ (
    .A(execution_unit_0.mab_lsb ),
    .Y(_01039_)
  );
  INVX1 _07341_ (
    .A(dbg_0.UNUSED_eu_mab_0_ ),
    .Y(_01040_)
  );
  INVX1 _07342_ (
    .A(execution_unit_0.mdb_in_buf_8_ ),
    .Y(_01041_)
  );
  INVX1 _07343_ (
    .A(execution_unit_0.mdb_in_buf_9_ ),
    .Y(_01042_)
  );
  INVX1 _07344_ (
    .A(execution_unit_0.mdb_in_buf_10_ ),
    .Y(_01043_)
  );
  INVX1 _07345_ (
    .A(execution_unit_0.mdb_in_buf_11_ ),
    .Y(_01044_)
  );
  INVX1 _07346_ (
    .A(execution_unit_0.mdb_in_buf_12_ ),
    .Y(_01045_)
  );
  INVX1 _07347_ (
    .A(execution_unit_0.mdb_in_buf_13_ ),
    .Y(_01046_)
  );
  INVX1 _07348_ (
    .A(execution_unit_0.mdb_in_buf_14_ ),
    .Y(_01047_)
  );
  INVX1 _07349_ (
    .A(execution_unit_0.mdb_in_buf_15_ ),
    .Y(_01048_)
  );
  INVX1 _07350_ (
    .A(dbg_0.dbg_reg_din_0_ ),
    .Y(_01049_)
  );
  INVX1 _07351_ (
    .A(dbg_0.dbg_reg_din_1_ ),
    .Y(_01050_)
  );
  INVX1 _07352_ (
    .A(dbg_0.dbg_reg_din_2_ ),
    .Y(_01051_)
  );
  INVX1 _07353_ (
    .A(dbg_0.dbg_reg_din_3_ ),
    .Y(_01052_)
  );
  INVX1 _07354_ (
    .A(dbg_0.dbg_reg_din_4_ ),
    .Y(_01053_)
  );
  INVX1 _07355_ (
    .A(dbg_0.dbg_reg_din_5_ ),
    .Y(_01054_)
  );
  INVX1 _07356_ (
    .A(dbg_0.dbg_reg_din_6_ ),
    .Y(_01055_)
  );
  INVX1 _07357_ (
    .A(dbg_0.dbg_reg_din_7_ ),
    .Y(_01056_)
  );
  INVX1 _07358_ (
    .A(dbg_0.dbg_reg_din_8_ ),
    .Y(_01057_)
  );
  INVX1 _07359_ (
    .A(dbg_0.dbg_reg_din_9_ ),
    .Y(_01058_)
  );
  INVX1 _07360_ (
    .A(dbg_0.dbg_reg_din_10_ ),
    .Y(_01059_)
  );
  INVX1 _07361_ (
    .A(dbg_0.dbg_reg_din_11_ ),
    .Y(_01060_)
  );
  INVX1 _07362_ (
    .A(dbg_0.dbg_reg_din_12_ ),
    .Y(_01061_)
  );
  INVX1 _07363_ (
    .A(dbg_0.dbg_reg_din_13_ ),
    .Y(_01062_)
  );
  INVX1 _07364_ (
    .A(dbg_0.dbg_reg_din_14_ ),
    .Y(_01063_)
  );
  INVX1 _07365_ (
    .A(dbg_0.dbg_reg_din_15_ ),
    .Y(_01064_)
  );
  INVX1 _07366_ (
    .A(cpu_halt_st),
    .Y(_01065_)
  );
  INVX1 _07367_ (
    .A(dbg_0.dbg_reg_wr ),
    .Y(_01066_)
  );
  INVX1 _07368_ (
    .A(_00162_),
    .Y(_01025_)
  );
  AND2X1 _07369_ (
    .A(_01027_),
    .B(e_state_3_),
    .Y(_01067_)
  );
  AND2X1 _07370_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .Y(_01068_)
  );
  NAND3X1 _07371_ (
    .A(_01027_),
    .B(e_state_3_),
    .C(_01068_),
    .Y(_01069_)
  );
  INVX1 _07372_ (
    .A(_01069_),
    .Y(execution_unit_0.alu_0.exec_cycle )
  );
  NOR2X1 _07373_ (
    .A(_01027_),
    .B(e_state_3_),
    .Y(_01070_)
  );
  NAND2X1 _07374_ (
    .A(e_state_1_),
    .B(_01070_),
    .Y(_01071_)
  );
  AND2X1 _07375_ (
    .A(_01026_),
    .B(e_state_1_),
    .Y(_01072_)
  );
  NAND2X1 _07376_ (
    .A(_01070_),
    .B(_01072_),
    .Y(_01073_)
  );
  INVX1 _07377_ (
    .A(_01073_),
    .Y(_01007_)
  );
  NOR2X1 _07378_ (
    .A(e_state_2_),
    .B(e_state_3_),
    .Y(_01074_)
  );
  NAND2X1 _07379_ (
    .A(_01026_),
    .B(_01074_),
    .Y(_01075_)
  );
  NOR2X1 _07380_ (
    .A(e_state_1_),
    .B(_01075_),
    .Y(execution_unit_0.reg_sr_clr )
  );
  NOR2X1 _07381_ (
    .A(_01026_),
    .B(e_state_1_),
    .Y(_01076_)
  );
  AND2X1 _07382_ (
    .A(_01067_),
    .B(_01076_),
    .Y(_01077_)
  );
  NAND2X1 _07383_ (
    .A(_01067_),
    .B(_01076_),
    .Y(_01078_)
  );
  OAI21X1 _07384_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(_01069_),
    .C(_01075_),
    .Y(_01079_)
  );
  MUX2X1 _07385_ (
    .A(execution_unit_0.alu_0.alu_out_0_ ),
    .B(eu_mdb_out_0_),
    .S(_01079_),
    .Y(_01080_)
  );
  NAND2X1 _07386_ (
    .A(UNUSED_fe_mab_0),
    .B(_01077_),
    .Y(_01081_)
  );
  OAI21X1 _07387_ (
    .A(_01077_),
    .B(_01080_),
    .C(_01081_),
    .Y(_01009_)
  );
  MUX2X1 _07388_ (
    .A(execution_unit_0.alu_0.alu_out_1_ ),
    .B(eu_mdb_out_1_),
    .S(_01079_),
    .Y(_01082_)
  );
  NAND2X1 _07389_ (
    .A(execution_unit_0.pc_nxt_1_ ),
    .B(_01077_),
    .Y(_01083_)
  );
  OAI21X1 _07390_ (
    .A(_01077_),
    .B(_01082_),
    .C(_01083_),
    .Y(_01016_)
  );
  MUX2X1 _07391_ (
    .A(execution_unit_0.alu_0.alu_out_2_ ),
    .B(eu_mdb_out_2_),
    .S(_01079_),
    .Y(_01084_)
  );
  NAND2X1 _07392_ (
    .A(execution_unit_0.pc_nxt_2_ ),
    .B(_01077_),
    .Y(_01085_)
  );
  OAI21X1 _07393_ (
    .A(_01077_),
    .B(_01084_),
    .C(_01085_),
    .Y(_01017_)
  );
  MUX2X1 _07394_ (
    .A(execution_unit_0.alu_0.alu_out_3_ ),
    .B(eu_mdb_out_3_),
    .S(_01079_),
    .Y(_01086_)
  );
  NAND2X1 _07395_ (
    .A(execution_unit_0.pc_nxt_3_ ),
    .B(_01077_),
    .Y(_01087_)
  );
  OAI21X1 _07396_ (
    .A(_01077_),
    .B(_01086_),
    .C(_01087_),
    .Y(_01018_)
  );
  MUX2X1 _07397_ (
    .A(execution_unit_0.alu_0.alu_out_4_ ),
    .B(eu_mdb_out_4_),
    .S(_01079_),
    .Y(_01088_)
  );
  NAND2X1 _07398_ (
    .A(execution_unit_0.pc_nxt_4_ ),
    .B(_01077_),
    .Y(_01089_)
  );
  OAI21X1 _07399_ (
    .A(_01077_),
    .B(_01088_),
    .C(_01089_),
    .Y(_01019_)
  );
  MUX2X1 _07400_ (
    .A(execution_unit_0.alu_0.alu_out_5_ ),
    .B(eu_mdb_out_5_),
    .S(_01079_),
    .Y(_01090_)
  );
  NAND2X1 _07401_ (
    .A(execution_unit_0.pc_nxt_5_ ),
    .B(_01077_),
    .Y(_01091_)
  );
  OAI21X1 _07402_ (
    .A(_01077_),
    .B(_01090_),
    .C(_01091_),
    .Y(_01020_)
  );
  MUX2X1 _07403_ (
    .A(execution_unit_0.alu_0.alu_out_6_ ),
    .B(eu_mdb_out_6_),
    .S(_01079_),
    .Y(_01092_)
  );
  NAND2X1 _07404_ (
    .A(execution_unit_0.pc_nxt_6_ ),
    .B(_01077_),
    .Y(_01093_)
  );
  OAI21X1 _07405_ (
    .A(_01077_),
    .B(_01092_),
    .C(_01093_),
    .Y(_01021_)
  );
  MUX2X1 _07406_ (
    .A(execution_unit_0.alu_0.alu_out_7_ ),
    .B(eu_mdb_out_7_),
    .S(_01079_),
    .Y(_01094_)
  );
  NAND2X1 _07407_ (
    .A(execution_unit_0.pc_nxt_7_ ),
    .B(_01077_),
    .Y(_01095_)
  );
  OAI21X1 _07408_ (
    .A(_01077_),
    .B(_01094_),
    .C(_01095_),
    .Y(_01022_)
  );
  MUX2X1 _07409_ (
    .A(execution_unit_0.alu_0.alu_out_8_ ),
    .B(execution_unit_0.mdb_out_nxt_8_ ),
    .S(_01079_),
    .Y(_01096_)
  );
  NAND2X1 _07410_ (
    .A(execution_unit_0.pc_nxt_8_ ),
    .B(_01077_),
    .Y(_01097_)
  );
  OAI21X1 _07411_ (
    .A(_01077_),
    .B(_01096_),
    .C(_01097_),
    .Y(_01023_)
  );
  MUX2X1 _07412_ (
    .A(execution_unit_0.alu_0.alu_out_9_ ),
    .B(execution_unit_0.mdb_out_nxt_9_ ),
    .S(_01079_),
    .Y(_01098_)
  );
  NAND2X1 _07413_ (
    .A(execution_unit_0.pc_nxt_9_ ),
    .B(_01077_),
    .Y(_01099_)
  );
  OAI21X1 _07414_ (
    .A(_01077_),
    .B(_01098_),
    .C(_01099_),
    .Y(_01024_)
  );
  MUX2X1 _07415_ (
    .A(execution_unit_0.alu_0.alu_out_10_ ),
    .B(execution_unit_0.mdb_out_nxt_10_ ),
    .S(_01079_),
    .Y(_01100_)
  );
  NAND2X1 _07416_ (
    .A(execution_unit_0.pc_nxt_10_ ),
    .B(_01077_),
    .Y(_01101_)
  );
  OAI21X1 _07417_ (
    .A(_01077_),
    .B(_01100_),
    .C(_01101_),
    .Y(_01010_)
  );
  MUX2X1 _07418_ (
    .A(execution_unit_0.alu_0.alu_out_11_ ),
    .B(execution_unit_0.mdb_out_nxt_11_ ),
    .S(_01079_),
    .Y(_01102_)
  );
  NAND2X1 _07419_ (
    .A(execution_unit_0.pc_nxt_11_ ),
    .B(_01077_),
    .Y(_01103_)
  );
  OAI21X1 _07420_ (
    .A(_01077_),
    .B(_01102_),
    .C(_01103_),
    .Y(_01011_)
  );
  MUX2X1 _07421_ (
    .A(execution_unit_0.alu_0.alu_out_12_ ),
    .B(execution_unit_0.mdb_out_nxt_12_ ),
    .S(_01079_),
    .Y(_01104_)
  );
  NAND2X1 _07422_ (
    .A(execution_unit_0.pc_nxt_12_ ),
    .B(_01077_),
    .Y(_01105_)
  );
  OAI21X1 _07423_ (
    .A(_01077_),
    .B(_01104_),
    .C(_01105_),
    .Y(_01012_)
  );
  MUX2X1 _07424_ (
    .A(execution_unit_0.alu_0.alu_out_13_ ),
    .B(execution_unit_0.mdb_out_nxt_13_ ),
    .S(_01079_),
    .Y(_01106_)
  );
  NAND2X1 _07425_ (
    .A(execution_unit_0.pc_nxt_13_ ),
    .B(_01077_),
    .Y(_01107_)
  );
  OAI21X1 _07426_ (
    .A(_01077_),
    .B(_01106_),
    .C(_01107_),
    .Y(_01013_)
  );
  MUX2X1 _07427_ (
    .A(execution_unit_0.alu_0.alu_out_14_ ),
    .B(execution_unit_0.mdb_out_nxt_14_ ),
    .S(_01079_),
    .Y(_01108_)
  );
  NAND2X1 _07428_ (
    .A(execution_unit_0.pc_nxt_14_ ),
    .B(_01077_),
    .Y(_01109_)
  );
  OAI21X1 _07429_ (
    .A(_01077_),
    .B(_01108_),
    .C(_01109_),
    .Y(_01014_)
  );
  MUX2X1 _07430_ (
    .A(execution_unit_0.alu_0.alu_out_15_ ),
    .B(execution_unit_0.mdb_out_nxt_15_ ),
    .S(_01079_),
    .Y(_01110_)
  );
  NAND2X1 _07431_ (
    .A(execution_unit_0.pc_nxt_15_ ),
    .B(_01077_),
    .Y(_01111_)
  );
  OAI21X1 _07432_ (
    .A(_01077_),
    .B(_01110_),
    .C(_01111_),
    .Y(_01015_)
  );
  NAND2X1 _07433_ (
    .A(e_state_0_),
    .B(_01074_),
    .Y(_01112_)
  );
  NOR2X1 _07434_ (
    .A(execution_unit_0.inst_irq_rst ),
    .B(_01112_),
    .Y(_01113_)
  );
  NAND2X1 _07435_ (
    .A(_01068_),
    .B(_01070_),
    .Y(_01114_)
  );
  NAND2X1 _07436_ (
    .A(_01067_),
    .B(_01072_),
    .Y(_01115_)
  );
  NAND3X1 _07437_ (
    .A(_01037_),
    .B(_01067_),
    .C(_01072_),
    .Y(_01116_)
  );
  OAI21X1 _07438_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01115_),
    .C(_01114_),
    .Y(_01117_)
  );
  OAI21X1 _07439_ (
    .A(_01113_),
    .B(_01117_),
    .C(_01038_),
    .Y(_01118_)
  );
  NOR2X1 _07440_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(execution_unit_0.inst_mov ),
    .Y(_01119_)
  );
  NAND2X1 _07441_ (
    .A(_01077_),
    .B(_01119_),
    .Y(_01120_)
  );
  OAI21X1 _07442_ (
    .A(execution_unit_0.inst_as_5_ ),
    .B(_01073_),
    .C(_01120_),
    .Y(_01121_)
  );
  AOI21X1 _07443_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(execution_unit_0.alu_0.exec_cycle ),
    .C(_01121_),
    .Y(_01122_)
  );
  NAND2X1 _07444_ (
    .A(_01118_),
    .B(_01122_),
    .Y(dbg_0.UNUSED_eu_mb_en )
  );
  MUX2X1 _07445_ (
    .A(_01040_),
    .B(_01039_),
    .S(dbg_0.UNUSED_eu_mb_en ),
    .Y(_00990_)
  );
  NAND2X1 _07446_ (
    .A(execution_unit_0.mab_lsb ),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01123_)
  );
  MUX2X1 _07447_ (
    .A(eu_mdb_in_0_),
    .B(eu_mdb_in_8_),
    .S(_01123_),
    .Y(_01124_)
  );
  NOR2X1 _07448_ (
    .A(execution_unit_0.mdb_in_buf_0_ ),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01125_)
  );
  AOI21X1 _07449_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01124_),
    .C(_01125_),
    .Y(_00991_)
  );
  MUX2X1 _07450_ (
    .A(eu_mdb_in_1_),
    .B(eu_mdb_in_9_),
    .S(_01123_),
    .Y(_01126_)
  );
  NOR2X1 _07451_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(execution_unit_0.mdb_in_buf_1_ ),
    .Y(_01127_)
  );
  AOI21X1 _07452_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01126_),
    .C(_01127_),
    .Y(_00998_)
  );
  MUX2X1 _07453_ (
    .A(eu_mdb_in_2_),
    .B(eu_mdb_in_10_),
    .S(_01123_),
    .Y(_01128_)
  );
  NOR2X1 _07454_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(execution_unit_0.mdb_in_buf_2_ ),
    .Y(_01129_)
  );
  AOI21X1 _07455_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01128_),
    .C(_01129_),
    .Y(_00999_)
  );
  MUX2X1 _07456_ (
    .A(eu_mdb_in_3_),
    .B(eu_mdb_in_11_),
    .S(_01123_),
    .Y(_01130_)
  );
  NOR2X1 _07457_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(execution_unit_0.mdb_in_buf_3_ ),
    .Y(_01131_)
  );
  AOI21X1 _07458_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01130_),
    .C(_01131_),
    .Y(_01000_)
  );
  MUX2X1 _07459_ (
    .A(eu_mdb_in_4_),
    .B(eu_mdb_in_12_),
    .S(_01123_),
    .Y(_01132_)
  );
  NOR2X1 _07460_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(execution_unit_0.mdb_in_buf_4_ ),
    .Y(_01133_)
  );
  AOI21X1 _07461_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01132_),
    .C(_01133_),
    .Y(_01001_)
  );
  MUX2X1 _07462_ (
    .A(eu_mdb_in_5_),
    .B(eu_mdb_in_13_),
    .S(_01123_),
    .Y(_01134_)
  );
  NOR2X1 _07463_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(execution_unit_0.mdb_in_buf_5_ ),
    .Y(_01135_)
  );
  AOI21X1 _07464_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01134_),
    .C(_01135_),
    .Y(_01002_)
  );
  MUX2X1 _07465_ (
    .A(eu_mdb_in_6_),
    .B(eu_mdb_in_14_),
    .S(_01123_),
    .Y(_01136_)
  );
  NOR2X1 _07466_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(execution_unit_0.mdb_in_buf_6_ ),
    .Y(_01137_)
  );
  AOI21X1 _07467_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01136_),
    .C(_01137_),
    .Y(_01003_)
  );
  MUX2X1 _07468_ (
    .A(eu_mdb_in_7_),
    .B(eu_mdb_in_15_),
    .S(_01123_),
    .Y(_01138_)
  );
  NOR2X1 _07469_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(execution_unit_0.mdb_in_buf_7_ ),
    .Y(_01139_)
  );
  AOI21X1 _07470_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01138_),
    .C(_01139_),
    .Y(_01004_)
  );
  NAND2X1 _07471_ (
    .A(eu_mdb_in_8_),
    .B(execution_unit_0.mdb_in_buf_en ),
    .Y(_01140_)
  );
  OAI21X1 _07472_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01041_),
    .C(_01140_),
    .Y(_01005_)
  );
  NAND2X1 _07473_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(eu_mdb_in_9_),
    .Y(_01141_)
  );
  OAI21X1 _07474_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01042_),
    .C(_01141_),
    .Y(_01006_)
  );
  NAND2X1 _07475_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(eu_mdb_in_10_),
    .Y(_01142_)
  );
  OAI21X1 _07476_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01043_),
    .C(_01142_),
    .Y(_00992_)
  );
  NAND2X1 _07477_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(eu_mdb_in_11_),
    .Y(_01143_)
  );
  OAI21X1 _07478_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01044_),
    .C(_01143_),
    .Y(_00993_)
  );
  NAND2X1 _07479_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(eu_mdb_in_12_),
    .Y(_01144_)
  );
  OAI21X1 _07480_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01045_),
    .C(_01144_),
    .Y(_00994_)
  );
  NAND2X1 _07481_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(eu_mdb_in_13_),
    .Y(_01145_)
  );
  OAI21X1 _07482_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01046_),
    .C(_01145_),
    .Y(_00995_)
  );
  NAND2X1 _07483_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(eu_mdb_in_14_),
    .Y(_01146_)
  );
  OAI21X1 _07484_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01047_),
    .C(_01146_),
    .Y(_00996_)
  );
  NAND2X1 _07485_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(eu_mdb_in_15_),
    .Y(_01147_)
  );
  OAI21X1 _07486_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(_01048_),
    .C(_01147_),
    .Y(_00997_)
  );
  OAI21X1 _07487_ (
    .A(execution_unit_0.mdb_in_buf_en ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01069_),
    .Y(_01148_)
  );
  INVX1 _07488_ (
    .A(_01148_),
    .Y(_01008_)
  );
  NOR2X1 _07489_ (
    .A(_01037_),
    .B(_01078_),
    .Y(execution_unit_0.reg_sr_wr )
  );
  NOR2X1 _07490_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .Y(_01149_)
  );
  OR2X1 _07491_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .Y(_01150_)
  );
  NOR3X1 _07492_ (
    .A(_01026_),
    .B(e_state_1_),
    .C(_01149_),
    .Y(_01151_)
  );
  NAND2X1 _07493_ (
    .A(_01067_),
    .B(_01151_),
    .Y(_01152_)
  );
  NAND3X1 _07494_ (
    .A(execution_unit_0.inst_as_1_ ),
    .B(_01070_),
    .C(_01151_),
    .Y(_01153_)
  );
  OAI21X1 _07495_ (
    .A(_01078_),
    .B(_01149_),
    .C(_01153_),
    .Y(_01154_)
  );
  AOI21X1 _07496_ (
    .A(e_state_0_),
    .B(_01074_),
    .C(_01154_),
    .Y(_01155_)
  );
  NOR2X1 _07497_ (
    .A(execution_unit_0.inst_as_3_ ),
    .B(execution_unit_0.inst_as_2_ ),
    .Y(_01156_)
  );
  OR2X1 _07498_ (
    .A(execution_unit_0.inst_as_6_ ),
    .B(execution_unit_0.inst_as_1_ ),
    .Y(_01157_)
  );
  NOR2X1 _07499_ (
    .A(execution_unit_0.inst_as_4_ ),
    .B(_01157_),
    .Y(_01158_)
  );
  AOI21X1 _07500_ (
    .A(_01156_),
    .B(_01158_),
    .C(_01069_),
    .Y(_01159_)
  );
  NOR2X1 _07501_ (
    .A(execution_unit_0.reg_sr_wr ),
    .B(_01159_),
    .Y(_01160_)
  );
  AOI21X1 _07502_ (
    .A(_01078_),
    .B(_01116_),
    .C(_01150_),
    .Y(_01161_)
  );
  NOR2X1 _07503_ (
    .A(execution_unit_0.inst_type_1_ ),
    .B(execution_unit_0.inst_as_7_ ),
    .Y(_01162_)
  );
  NOR2X1 _07504_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(execution_unit_0.inst_as_5_ ),
    .Y(_01163_)
  );
  AOI21X1 _07505_ (
    .A(_01162_),
    .B(_01163_),
    .C(_01069_),
    .Y(_01164_)
  );
  AOI22X1 _07506_ (
    .A(execution_unit_0.inst_dext_0_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_0_ ),
    .Y(_01165_)
  );
  NOR2X1 _07507_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01124_),
    .Y(_01166_)
  );
  AOI21X1 _07508_ (
    .A(execution_unit_0.mdb_in_buf_0_ ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01166_),
    .Y(_01167_)
  );
  MUX2X1 _07509_ (
    .A(_01165_),
    .B(_01167_),
    .S(_01160_),
    .Y(_01168_)
  );
  NOR2X1 _07510_ (
    .A(execution_unit_0.inst_type_1_ ),
    .B(_01069_),
    .Y(_01169_)
  );
  AOI22X1 _07511_ (
    .A(_01026_),
    .B(_01074_),
    .C(_01169_),
    .D(execution_unit_0.inst_as_0_ ),
    .Y(_01170_)
  );
  OAI21X1 _07512_ (
    .A(execution_unit_0.inst_as_6_ ),
    .B(_01071_),
    .C(_01170_),
    .Y(_01171_)
  );
  MUX2X1 _07513_ (
    .A(_01168_),
    .B(dbg_0.dbg_reg_din_0_ ),
    .S(_01155_),
    .Y(_01172_)
  );
  NAND2X1 _07514_ (
    .A(execution_unit_0.reg_src_0_ ),
    .B(_01171_),
    .Y(_01173_)
  );
  OAI21X1 _07515_ (
    .A(_01171_),
    .B(_01172_),
    .C(_01173_),
    .Y(execution_unit_0.alu_0.alu_swpb_8_ )
  );
  AOI22X1 _07516_ (
    .A(execution_unit_0.inst_dext_1_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_1_ ),
    .Y(_01174_)
  );
  NOR2X1 _07517_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01126_),
    .Y(_01175_)
  );
  AOI21X1 _07518_ (
    .A(execution_unit_0.mdb_in_buf_1_ ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01175_),
    .Y(_01176_)
  );
  MUX2X1 _07519_ (
    .A(_01174_),
    .B(_01176_),
    .S(_01160_),
    .Y(_01177_)
  );
  MUX2X1 _07520_ (
    .A(_01177_),
    .B(dbg_0.dbg_reg_din_1_ ),
    .S(_01155_),
    .Y(_01178_)
  );
  NAND2X1 _07521_ (
    .A(execution_unit_0.reg_src_1_ ),
    .B(_01171_),
    .Y(_01179_)
  );
  OAI21X1 _07522_ (
    .A(_01171_),
    .B(_01178_),
    .C(_01179_),
    .Y(execution_unit_0.alu_0.alu_shift_0_ )
  );
  AOI22X1 _07523_ (
    .A(execution_unit_0.inst_dext_2_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_2_ ),
    .Y(_01180_)
  );
  NOR2X1 _07524_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01128_),
    .Y(_01181_)
  );
  AOI21X1 _07525_ (
    .A(execution_unit_0.mdb_in_buf_2_ ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01181_),
    .Y(_01182_)
  );
  MUX2X1 _07526_ (
    .A(_01180_),
    .B(_01182_),
    .S(_01160_),
    .Y(_01183_)
  );
  MUX2X1 _07527_ (
    .A(_01183_),
    .B(dbg_0.dbg_reg_din_2_ ),
    .S(_01155_),
    .Y(_01184_)
  );
  NAND2X1 _07528_ (
    .A(execution_unit_0.reg_src_2_ ),
    .B(_01171_),
    .Y(_01185_)
  );
  OAI21X1 _07529_ (
    .A(_01171_),
    .B(_01184_),
    .C(_01185_),
    .Y(execution_unit_0.alu_0.alu_shift_1_ )
  );
  AOI22X1 _07530_ (
    .A(execution_unit_0.inst_dext_3_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_3_ ),
    .Y(_01186_)
  );
  NOR2X1 _07531_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01130_),
    .Y(_01187_)
  );
  AOI21X1 _07532_ (
    .A(execution_unit_0.mdb_in_buf_3_ ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01187_),
    .Y(_01188_)
  );
  MUX2X1 _07533_ (
    .A(_01186_),
    .B(_01188_),
    .S(_01160_),
    .Y(_01189_)
  );
  MUX2X1 _07534_ (
    .A(_01189_),
    .B(dbg_0.dbg_reg_din_3_ ),
    .S(_01155_),
    .Y(_01190_)
  );
  NAND2X1 _07535_ (
    .A(execution_unit_0.reg_src_3_ ),
    .B(_01171_),
    .Y(_01191_)
  );
  OAI21X1 _07536_ (
    .A(_01171_),
    .B(_01190_),
    .C(_01191_),
    .Y(execution_unit_0.alu_0.alu_shift_2_ )
  );
  AOI22X1 _07537_ (
    .A(execution_unit_0.inst_dext_4_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_4_ ),
    .Y(_01192_)
  );
  NOR2X1 _07538_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01132_),
    .Y(_01193_)
  );
  AOI21X1 _07539_ (
    .A(execution_unit_0.mdb_in_buf_4_ ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01193_),
    .Y(_01194_)
  );
  MUX2X1 _07540_ (
    .A(_01192_),
    .B(_01194_),
    .S(_01160_),
    .Y(_01195_)
  );
  MUX2X1 _07541_ (
    .A(_01195_),
    .B(dbg_0.dbg_reg_din_4_ ),
    .S(_01155_),
    .Y(_01196_)
  );
  NAND2X1 _07542_ (
    .A(execution_unit_0.reg_src_4_ ),
    .B(_01171_),
    .Y(_01197_)
  );
  OAI21X1 _07543_ (
    .A(_01171_),
    .B(_01196_),
    .C(_01197_),
    .Y(execution_unit_0.alu_0.alu_shift_3_ )
  );
  AOI22X1 _07544_ (
    .A(execution_unit_0.inst_dext_5_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_5_ ),
    .Y(_01198_)
  );
  NOR2X1 _07545_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01134_),
    .Y(_01199_)
  );
  AOI21X1 _07546_ (
    .A(execution_unit_0.mdb_in_buf_5_ ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01199_),
    .Y(_01200_)
  );
  MUX2X1 _07547_ (
    .A(_01198_),
    .B(_01200_),
    .S(_01160_),
    .Y(_01201_)
  );
  MUX2X1 _07548_ (
    .A(_01201_),
    .B(dbg_0.dbg_reg_din_5_ ),
    .S(_01155_),
    .Y(_01202_)
  );
  NAND2X1 _07549_ (
    .A(execution_unit_0.reg_src_5_ ),
    .B(_01171_),
    .Y(_01203_)
  );
  OAI21X1 _07550_ (
    .A(_01171_),
    .B(_01202_),
    .C(_01203_),
    .Y(execution_unit_0.alu_0.alu_shift_4_ )
  );
  AOI22X1 _07551_ (
    .A(execution_unit_0.inst_dext_6_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_6_ ),
    .Y(_01204_)
  );
  NOR2X1 _07552_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01136_),
    .Y(_01205_)
  );
  AOI21X1 _07553_ (
    .A(execution_unit_0.mdb_in_buf_6_ ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01205_),
    .Y(_01206_)
  );
  MUX2X1 _07554_ (
    .A(_01204_),
    .B(_01206_),
    .S(_01160_),
    .Y(_01207_)
  );
  MUX2X1 _07555_ (
    .A(_01207_),
    .B(dbg_0.dbg_reg_din_6_ ),
    .S(_01155_),
    .Y(_01208_)
  );
  NAND2X1 _07556_ (
    .A(execution_unit_0.reg_src_6_ ),
    .B(_01171_),
    .Y(_01209_)
  );
  OAI21X1 _07557_ (
    .A(_01171_),
    .B(_01208_),
    .C(_01209_),
    .Y(execution_unit_0.alu_0.alu_shift_5_ )
  );
  AOI22X1 _07558_ (
    .A(execution_unit_0.inst_dext_7_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_7_ ),
    .Y(_01210_)
  );
  NOR2X1 _07559_ (
    .A(execution_unit_0.mdb_in_buf_valid ),
    .B(_01138_),
    .Y(_01211_)
  );
  AOI21X1 _07560_ (
    .A(execution_unit_0.mdb_in_buf_7_ ),
    .B(execution_unit_0.mdb_in_buf_valid ),
    .C(_01211_),
    .Y(_01212_)
  );
  MUX2X1 _07561_ (
    .A(_01210_),
    .B(_01212_),
    .S(_01160_),
    .Y(_01213_)
  );
  MUX2X1 _07562_ (
    .A(_01213_),
    .B(dbg_0.dbg_reg_din_7_ ),
    .S(_01155_),
    .Y(_01214_)
  );
  NAND2X1 _07563_ (
    .A(execution_unit_0.reg_src_7_ ),
    .B(_01171_),
    .Y(_01215_)
  );
  OAI21X1 _07564_ (
    .A(_01171_),
    .B(_01214_),
    .C(_01215_),
    .Y(execution_unit_0.alu_0.alu_shift_6_ )
  );
  AOI22X1 _07565_ (
    .A(execution_unit_0.inst_dext_8_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_8_ ),
    .Y(_01216_)
  );
  MUX2X1 _07566_ (
    .A(execution_unit_0.mdb_in_buf_8_ ),
    .B(eu_mdb_in_8_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01217_)
  );
  MUX2X1 _07567_ (
    .A(_01216_),
    .B(_01217_),
    .S(_01160_),
    .Y(_01218_)
  );
  MUX2X1 _07568_ (
    .A(_01218_),
    .B(dbg_0.dbg_reg_din_8_ ),
    .S(_01155_),
    .Y(_01219_)
  );
  NAND2X1 _07569_ (
    .A(execution_unit_0.reg_src_8_ ),
    .B(_01171_),
    .Y(_01220_)
  );
  OAI21X1 _07570_ (
    .A(_01171_),
    .B(_01219_),
    .C(_01220_),
    .Y(execution_unit_0.alu_0.alu_swpb_0_ )
  );
  AOI22X1 _07571_ (
    .A(execution_unit_0.inst_dext_9_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_9_ ),
    .Y(_01221_)
  );
  MUX2X1 _07572_ (
    .A(execution_unit_0.mdb_in_buf_9_ ),
    .B(eu_mdb_in_9_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01222_)
  );
  MUX2X1 _07573_ (
    .A(_01221_),
    .B(_01222_),
    .S(_01160_),
    .Y(_01223_)
  );
  MUX2X1 _07574_ (
    .A(_01223_),
    .B(dbg_0.dbg_reg_din_9_ ),
    .S(_01155_),
    .Y(_01224_)
  );
  NAND2X1 _07575_ (
    .A(execution_unit_0.reg_src_9_ ),
    .B(_01171_),
    .Y(_01225_)
  );
  OAI21X1 _07576_ (
    .A(_01171_),
    .B(_01224_),
    .C(_01225_),
    .Y(execution_unit_0.alu_0.alu_shift_8_ )
  );
  AOI22X1 _07577_ (
    .A(execution_unit_0.inst_dext_10_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_10_ ),
    .Y(_01226_)
  );
  MUX2X1 _07578_ (
    .A(execution_unit_0.mdb_in_buf_10_ ),
    .B(eu_mdb_in_10_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01227_)
  );
  MUX2X1 _07579_ (
    .A(_01226_),
    .B(_01227_),
    .S(_01160_),
    .Y(_01228_)
  );
  MUX2X1 _07580_ (
    .A(_01228_),
    .B(dbg_0.dbg_reg_din_10_ ),
    .S(_01155_),
    .Y(_01229_)
  );
  NAND2X1 _07581_ (
    .A(execution_unit_0.reg_src_10_ ),
    .B(_01171_),
    .Y(_01230_)
  );
  OAI21X1 _07582_ (
    .A(_01171_),
    .B(_01229_),
    .C(_01230_),
    .Y(execution_unit_0.alu_0.alu_shift_9_ )
  );
  AOI22X1 _07583_ (
    .A(execution_unit_0.inst_dext_11_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_11_ ),
    .Y(_01231_)
  );
  MUX2X1 _07584_ (
    .A(execution_unit_0.mdb_in_buf_11_ ),
    .B(eu_mdb_in_11_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01232_)
  );
  MUX2X1 _07585_ (
    .A(_01231_),
    .B(_01232_),
    .S(_01160_),
    .Y(_01233_)
  );
  MUX2X1 _07586_ (
    .A(_01233_),
    .B(dbg_0.dbg_reg_din_11_ ),
    .S(_01155_),
    .Y(_01234_)
  );
  NAND2X1 _07587_ (
    .A(execution_unit_0.reg_src_11_ ),
    .B(_01171_),
    .Y(_01235_)
  );
  OAI21X1 _07588_ (
    .A(_01171_),
    .B(_01234_),
    .C(_01235_),
    .Y(execution_unit_0.alu_0.alu_shift_10_ )
  );
  AOI22X1 _07589_ (
    .A(execution_unit_0.inst_dext_12_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_12_ ),
    .Y(_01236_)
  );
  MUX2X1 _07590_ (
    .A(execution_unit_0.mdb_in_buf_12_ ),
    .B(eu_mdb_in_12_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01237_)
  );
  MUX2X1 _07591_ (
    .A(_01236_),
    .B(_01237_),
    .S(_01160_),
    .Y(_01238_)
  );
  MUX2X1 _07592_ (
    .A(_01238_),
    .B(dbg_0.dbg_reg_din_12_ ),
    .S(_01155_),
    .Y(_01239_)
  );
  NAND2X1 _07593_ (
    .A(execution_unit_0.reg_src_12_ ),
    .B(_01171_),
    .Y(_01240_)
  );
  OAI21X1 _07594_ (
    .A(_01171_),
    .B(_01239_),
    .C(_01240_),
    .Y(execution_unit_0.alu_0.alu_shift_11_ )
  );
  AOI22X1 _07595_ (
    .A(execution_unit_0.inst_dext_13_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_13_ ),
    .Y(_01241_)
  );
  MUX2X1 _07596_ (
    .A(execution_unit_0.mdb_in_buf_13_ ),
    .B(eu_mdb_in_13_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01242_)
  );
  MUX2X1 _07597_ (
    .A(_01241_),
    .B(_01242_),
    .S(_01160_),
    .Y(_01243_)
  );
  MUX2X1 _07598_ (
    .A(_01243_),
    .B(dbg_0.dbg_reg_din_13_ ),
    .S(_01155_),
    .Y(_01244_)
  );
  NAND2X1 _07599_ (
    .A(execution_unit_0.reg_src_13_ ),
    .B(_01171_),
    .Y(_01245_)
  );
  OAI21X1 _07600_ (
    .A(_01171_),
    .B(_01244_),
    .C(_01245_),
    .Y(execution_unit_0.alu_0.alu_shift_12_ )
  );
  AOI22X1 _07601_ (
    .A(execution_unit_0.inst_dext_14_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_14_ ),
    .Y(_01246_)
  );
  MUX2X1 _07602_ (
    .A(execution_unit_0.mdb_in_buf_14_ ),
    .B(eu_mdb_in_14_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01247_)
  );
  MUX2X1 _07603_ (
    .A(_01246_),
    .B(_01247_),
    .S(_01160_),
    .Y(_01248_)
  );
  MUX2X1 _07604_ (
    .A(_01248_),
    .B(dbg_0.dbg_reg_din_14_ ),
    .S(_01155_),
    .Y(_01249_)
  );
  NAND2X1 _07605_ (
    .A(execution_unit_0.reg_src_14_ ),
    .B(_01171_),
    .Y(_01250_)
  );
  OAI21X1 _07606_ (
    .A(_01171_),
    .B(_01249_),
    .C(_01250_),
    .Y(execution_unit_0.alu_0.alu_shift_13_ )
  );
  AOI22X1 _07607_ (
    .A(execution_unit_0.inst_dext_15_ ),
    .B(_01161_),
    .C(_01164_),
    .D(execution_unit_0.inst_sext_15_ ),
    .Y(_01251_)
  );
  MUX2X1 _07608_ (
    .A(execution_unit_0.mdb_in_buf_15_ ),
    .B(eu_mdb_in_15_),
    .S(execution_unit_0.mdb_in_buf_valid ),
    .Y(_01252_)
  );
  MUX2X1 _07609_ (
    .A(_01251_),
    .B(_01252_),
    .S(_01160_),
    .Y(_01253_)
  );
  MUX2X1 _07610_ (
    .A(_01253_),
    .B(dbg_0.dbg_reg_din_15_ ),
    .S(_01155_),
    .Y(_01254_)
  );
  NAND2X1 _07611_ (
    .A(execution_unit_0.reg_src_15_ ),
    .B(_01171_),
    .Y(_01255_)
  );
  OAI21X1 _07612_ (
    .A(_01171_),
    .B(_01254_),
    .C(_01255_),
    .Y(execution_unit_0.alu_0.alu_shift_14_ )
  );
  NOR2X1 _07613_ (
    .A(_00144_),
    .B(_01065_),
    .Y(_01256_)
  );
  OR2X1 _07614_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(execution_unit_0.inst_type_1_ ),
    .Y(_01257_)
  );
  NOR2X1 _07615_ (
    .A(execution_unit_0.inst_ad_0_ ),
    .B(_01257_),
    .Y(_01258_)
  );
  INVX1 _07616_ (
    .A(_01258_),
    .Y(_01259_)
  );
  NOR2X1 _07617_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01069_),
    .Y(_01260_)
  );
  OR2X1 _07618_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01069_),
    .Y(_01261_)
  );
  NAND3X1 _07619_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01067_),
    .C(_01072_),
    .Y(_01262_)
  );
  INVX1 _07620_ (
    .A(_01262_),
    .Y(_01263_)
  );
  AOI21X1 _07621_ (
    .A(_01258_),
    .B(_01260_),
    .C(_01263_),
    .Y(_01264_)
  );
  OAI21X1 _07622_ (
    .A(_01259_),
    .B(_01261_),
    .C(_01262_),
    .Y(_01265_)
  );
  NOR2X1 _07623_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01150_),
    .Y(_01266_)
  );
  NAND3X1 _07624_ (
    .A(_01067_),
    .B(_01076_),
    .C(_01266_),
    .Y(_01267_)
  );
  AOI21X1 _07625_ (
    .A(_01115_),
    .B(_01267_),
    .C(execution_unit_0.inst_ad_6_ ),
    .Y(_01268_)
  );
  AOI21X1 _07626_ (
    .A(_01259_),
    .B(_01260_),
    .C(_01268_),
    .Y(_01269_)
  );
  OAI21X1 _07627_ (
    .A(_01049_),
    .B(_01269_),
    .C(_01264_),
    .Y(_01270_)
  );
  NAND2X1 _07628_ (
    .A(_01124_),
    .B(_01265_),
    .Y(_01271_)
  );
  NAND2X1 _07629_ (
    .A(_01270_),
    .B(_01271_),
    .Y(_01272_)
  );
  NOR2X1 _07630_ (
    .A(_01071_),
    .B(_01158_),
    .Y(_01273_)
  );
  OR2X1 _07631_ (
    .A(_01071_),
    .B(_01158_),
    .Y(_01274_)
  );
  AOI21X1 _07632_ (
    .A(execution_unit_0.inst_sext_0_ ),
    .B(_01273_),
    .C(cpu_halt_st),
    .Y(_01275_)
  );
  AOI21X1 _07633_ (
    .A(_01272_),
    .B(_01275_),
    .C(_01256_),
    .Y(execution_unit_0.alu_0.op_dst_0_ )
  );
  NAND2X1 _07634_ (
    .A(cpu_halt_st),
    .B(_00151_),
    .Y(_01276_)
  );
  OAI21X1 _07635_ (
    .A(execution_unit_0.inst_as_3_ ),
    .B(execution_unit_0.inst_as_2_ ),
    .C(execution_unit_0.inst_src_1_ ),
    .Y(_01277_)
  );
  INVX1 _07636_ (
    .A(_01277_),
    .Y(_01278_)
  );
  OAI21X1 _07637_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .C(_01278_),
    .Y(_01279_)
  );
  OAI21X1 _07638_ (
    .A(_01073_),
    .B(_01279_),
    .C(_01153_),
    .Y(_01280_)
  );
  OAI21X1 _07639_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .C(_01074_),
    .Y(_01281_)
  );
  OAI21X1 _07640_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_01152_),
    .C(_01281_),
    .Y(_01282_)
  );
  NOR3X1 _07641_ (
    .A(_01265_),
    .B(_01280_),
    .C(_01282_),
    .Y(_01283_)
  );
  OAI21X1 _07642_ (
    .A(_01050_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01284_)
  );
  NAND2X1 _07643_ (
    .A(_01126_),
    .B(_01265_),
    .Y(_01285_)
  );
  AOI21X1 _07644_ (
    .A(_01284_),
    .B(_01285_),
    .C(_01273_),
    .Y(_01286_)
  );
  OAI21X1 _07645_ (
    .A(execution_unit_0.inst_sext_1_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01287_)
  );
  OAI21X1 _07646_ (
    .A(_01286_),
    .B(_01287_),
    .C(_01276_),
    .Y(execution_unit_0.alu_0.op_dst_1_ )
  );
  NAND2X1 _07647_ (
    .A(cpu_halt_st),
    .B(_00152_),
    .Y(_01288_)
  );
  OAI21X1 _07648_ (
    .A(_01051_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01289_)
  );
  NAND2X1 _07649_ (
    .A(_01128_),
    .B(_01265_),
    .Y(_01290_)
  );
  AOI21X1 _07650_ (
    .A(_01289_),
    .B(_01290_),
    .C(_01273_),
    .Y(_01291_)
  );
  OAI21X1 _07651_ (
    .A(execution_unit_0.inst_sext_2_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01292_)
  );
  OAI21X1 _07652_ (
    .A(_01291_),
    .B(_01292_),
    .C(_01288_),
    .Y(execution_unit_0.alu_0.op_dst_2_ )
  );
  NAND2X1 _07653_ (
    .A(cpu_halt_st),
    .B(_00153_),
    .Y(_01293_)
  );
  OAI21X1 _07654_ (
    .A(_01052_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01294_)
  );
  NAND2X1 _07655_ (
    .A(_01130_),
    .B(_01265_),
    .Y(_01295_)
  );
  AOI21X1 _07656_ (
    .A(_01294_),
    .B(_01295_),
    .C(_01273_),
    .Y(_01296_)
  );
  OAI21X1 _07657_ (
    .A(execution_unit_0.inst_sext_3_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01297_)
  );
  OAI21X1 _07658_ (
    .A(_01296_),
    .B(_01297_),
    .C(_01293_),
    .Y(execution_unit_0.alu_0.op_dst_3_ )
  );
  NAND2X1 _07659_ (
    .A(cpu_halt_st),
    .B(_00154_),
    .Y(_01298_)
  );
  OAI21X1 _07660_ (
    .A(_01053_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01299_)
  );
  NAND2X1 _07661_ (
    .A(_01132_),
    .B(_01265_),
    .Y(_01300_)
  );
  AOI21X1 _07662_ (
    .A(_01299_),
    .B(_01300_),
    .C(_01273_),
    .Y(_01301_)
  );
  OAI21X1 _07663_ (
    .A(execution_unit_0.inst_sext_4_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01302_)
  );
  OAI21X1 _07664_ (
    .A(_01301_),
    .B(_01302_),
    .C(_01298_),
    .Y(execution_unit_0.alu_0.op_dst_4_ )
  );
  NAND2X1 _07665_ (
    .A(cpu_halt_st),
    .B(_00155_),
    .Y(_01303_)
  );
  OAI21X1 _07666_ (
    .A(_01054_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01304_)
  );
  NAND2X1 _07667_ (
    .A(_01134_),
    .B(_01265_),
    .Y(_01305_)
  );
  AOI21X1 _07668_ (
    .A(_01304_),
    .B(_01305_),
    .C(_01273_),
    .Y(_01306_)
  );
  OAI21X1 _07669_ (
    .A(execution_unit_0.inst_sext_5_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01307_)
  );
  OAI21X1 _07670_ (
    .A(_01306_),
    .B(_01307_),
    .C(_01303_),
    .Y(execution_unit_0.alu_0.op_dst_5_ )
  );
  NAND2X1 _07671_ (
    .A(cpu_halt_st),
    .B(_00156_),
    .Y(_01308_)
  );
  OAI21X1 _07672_ (
    .A(_01055_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01309_)
  );
  NAND2X1 _07673_ (
    .A(_01136_),
    .B(_01265_),
    .Y(_01310_)
  );
  AOI21X1 _07674_ (
    .A(_01309_),
    .B(_01310_),
    .C(_01273_),
    .Y(_01311_)
  );
  OAI21X1 _07675_ (
    .A(execution_unit_0.inst_sext_6_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01312_)
  );
  OAI21X1 _07676_ (
    .A(_01311_),
    .B(_01312_),
    .C(_01308_),
    .Y(execution_unit_0.alu_0.op_dst_6_ )
  );
  NAND2X1 _07677_ (
    .A(cpu_halt_st),
    .B(_00157_),
    .Y(_01313_)
  );
  OAI21X1 _07678_ (
    .A(_01056_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01314_)
  );
  NAND2X1 _07679_ (
    .A(_01138_),
    .B(_01265_),
    .Y(_01315_)
  );
  AOI21X1 _07680_ (
    .A(_01314_),
    .B(_01315_),
    .C(_01273_),
    .Y(_01316_)
  );
  OAI21X1 _07681_ (
    .A(execution_unit_0.inst_sext_7_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01317_)
  );
  OAI21X1 _07682_ (
    .A(_01316_),
    .B(_01317_),
    .C(_01313_),
    .Y(execution_unit_0.alu_0.op_dst_7_ )
  );
  NAND2X1 _07683_ (
    .A(cpu_halt_st),
    .B(_00158_),
    .Y(_01318_)
  );
  OAI21X1 _07684_ (
    .A(_01057_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01319_)
  );
  OR2X1 _07685_ (
    .A(eu_mdb_in_8_),
    .B(_01264_),
    .Y(_01320_)
  );
  AOI21X1 _07686_ (
    .A(_01319_),
    .B(_01320_),
    .C(_01273_),
    .Y(_01321_)
  );
  OAI21X1 _07687_ (
    .A(execution_unit_0.inst_sext_8_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01322_)
  );
  OAI21X1 _07688_ (
    .A(_01321_),
    .B(_01322_),
    .C(_01318_),
    .Y(execution_unit_0.alu_0.op_dst_8_ )
  );
  NAND2X1 _07689_ (
    .A(cpu_halt_st),
    .B(_00159_),
    .Y(_01323_)
  );
  OAI21X1 _07690_ (
    .A(_01058_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01324_)
  );
  OR2X1 _07691_ (
    .A(eu_mdb_in_9_),
    .B(_01264_),
    .Y(_01325_)
  );
  AOI21X1 _07692_ (
    .A(_01324_),
    .B(_01325_),
    .C(_01273_),
    .Y(_01326_)
  );
  OAI21X1 _07693_ (
    .A(execution_unit_0.inst_sext_9_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01327_)
  );
  OAI21X1 _07694_ (
    .A(_01326_),
    .B(_01327_),
    .C(_01323_),
    .Y(execution_unit_0.alu_0.op_dst_9_ )
  );
  NAND2X1 _07695_ (
    .A(cpu_halt_st),
    .B(_00145_),
    .Y(_01328_)
  );
  OAI21X1 _07696_ (
    .A(_01059_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01329_)
  );
  OR2X1 _07697_ (
    .A(eu_mdb_in_10_),
    .B(_01264_),
    .Y(_01330_)
  );
  AOI21X1 _07698_ (
    .A(_01329_),
    .B(_01330_),
    .C(_01273_),
    .Y(_01331_)
  );
  OAI21X1 _07699_ (
    .A(execution_unit_0.inst_sext_10_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01332_)
  );
  OAI21X1 _07700_ (
    .A(_01331_),
    .B(_01332_),
    .C(_01328_),
    .Y(execution_unit_0.alu_0.op_dst_10_ )
  );
  NAND2X1 _07701_ (
    .A(cpu_halt_st),
    .B(_00146_),
    .Y(_01333_)
  );
  OAI21X1 _07702_ (
    .A(_01060_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01334_)
  );
  OR2X1 _07703_ (
    .A(eu_mdb_in_11_),
    .B(_01264_),
    .Y(_01335_)
  );
  AOI21X1 _07704_ (
    .A(_01334_),
    .B(_01335_),
    .C(_01273_),
    .Y(_01336_)
  );
  OAI21X1 _07705_ (
    .A(execution_unit_0.inst_sext_11_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01337_)
  );
  OAI21X1 _07706_ (
    .A(_01336_),
    .B(_01337_),
    .C(_01333_),
    .Y(execution_unit_0.alu_0.op_dst_11_ )
  );
  NAND2X1 _07707_ (
    .A(cpu_halt_st),
    .B(_00147_),
    .Y(_01338_)
  );
  OAI21X1 _07708_ (
    .A(_01061_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01339_)
  );
  OR2X1 _07709_ (
    .A(eu_mdb_in_12_),
    .B(_01264_),
    .Y(_01340_)
  );
  AOI21X1 _07710_ (
    .A(_01339_),
    .B(_01340_),
    .C(_01273_),
    .Y(_01341_)
  );
  OAI21X1 _07711_ (
    .A(execution_unit_0.inst_sext_12_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01342_)
  );
  OAI21X1 _07712_ (
    .A(_01341_),
    .B(_01342_),
    .C(_01338_),
    .Y(execution_unit_0.alu_0.op_dst_12_ )
  );
  NAND2X1 _07713_ (
    .A(cpu_halt_st),
    .B(_00148_),
    .Y(_01343_)
  );
  OAI21X1 _07714_ (
    .A(_01062_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01344_)
  );
  OR2X1 _07715_ (
    .A(eu_mdb_in_13_),
    .B(_01264_),
    .Y(_01345_)
  );
  AOI21X1 _07716_ (
    .A(_01344_),
    .B(_01345_),
    .C(_01273_),
    .Y(_01346_)
  );
  OAI21X1 _07717_ (
    .A(execution_unit_0.inst_sext_13_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01347_)
  );
  OAI21X1 _07718_ (
    .A(_01346_),
    .B(_01347_),
    .C(_01343_),
    .Y(execution_unit_0.alu_0.op_dst_13_ )
  );
  NAND2X1 _07719_ (
    .A(cpu_halt_st),
    .B(_00149_),
    .Y(_01348_)
  );
  OAI21X1 _07720_ (
    .A(_01063_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01349_)
  );
  OR2X1 _07721_ (
    .A(eu_mdb_in_14_),
    .B(_01264_),
    .Y(_01350_)
  );
  AOI21X1 _07722_ (
    .A(_01349_),
    .B(_01350_),
    .C(_01273_),
    .Y(_01351_)
  );
  OAI21X1 _07723_ (
    .A(execution_unit_0.inst_sext_14_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01352_)
  );
  OAI21X1 _07724_ (
    .A(_01351_),
    .B(_01352_),
    .C(_01348_),
    .Y(execution_unit_0.alu_0.op_dst_14_ )
  );
  NAND2X1 _07725_ (
    .A(cpu_halt_st),
    .B(_00150_),
    .Y(_01353_)
  );
  OAI21X1 _07726_ (
    .A(_01064_),
    .B(_01269_),
    .C(_01283_),
    .Y(_01354_)
  );
  OR2X1 _07727_ (
    .A(eu_mdb_in_15_),
    .B(_01264_),
    .Y(_01355_)
  );
  AOI21X1 _07728_ (
    .A(_01354_),
    .B(_01355_),
    .C(_01273_),
    .Y(_01356_)
  );
  OAI21X1 _07729_ (
    .A(execution_unit_0.inst_sext_15_ ),
    .B(_01274_),
    .C(_01065_),
    .Y(_01357_)
  );
  OAI21X1 _07730_ (
    .A(_01356_),
    .B(_01357_),
    .C(_01353_),
    .Y(execution_unit_0.alu_0.op_dst_15_ )
  );
  NAND2X1 _07731_ (
    .A(eu_mdb_out_0_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01358_)
  );
  OAI21X1 _07732_ (
    .A(_01029_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01358_),
    .Y(eu_mdb_out_8_)
  );
  NAND2X1 _07733_ (
    .A(eu_mdb_out_1_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01359_)
  );
  OAI21X1 _07734_ (
    .A(_01030_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01359_),
    .Y(eu_mdb_out_9_)
  );
  NAND2X1 _07735_ (
    .A(eu_mdb_out_2_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01360_)
  );
  OAI21X1 _07736_ (
    .A(_01031_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01360_),
    .Y(eu_mdb_out_10_)
  );
  NAND2X1 _07737_ (
    .A(eu_mdb_out_3_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01361_)
  );
  OAI21X1 _07738_ (
    .A(_01032_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01361_),
    .Y(eu_mdb_out_11_)
  );
  NAND2X1 _07739_ (
    .A(eu_mdb_out_4_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01362_)
  );
  OAI21X1 _07740_ (
    .A(_01033_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01362_),
    .Y(eu_mdb_out_12_)
  );
  NAND2X1 _07741_ (
    .A(eu_mdb_out_5_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01363_)
  );
  OAI21X1 _07742_ (
    .A(_01034_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01363_),
    .Y(eu_mdb_out_13_)
  );
  NAND2X1 _07743_ (
    .A(eu_mdb_out_6_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01364_)
  );
  OAI21X1 _07744_ (
    .A(_01035_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01364_),
    .Y(eu_mdb_out_14_)
  );
  NAND2X1 _07745_ (
    .A(eu_mdb_out_7_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01365_)
  );
  OAI21X1 _07746_ (
    .A(_01036_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01365_),
    .Y(eu_mdb_out_15_)
  );
  NAND3X1 _07747_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(execution_unit_0.inst_as_0_ ),
    .C(_01266_),
    .Y(_01366_)
  );
  NAND2X1 _07748_ (
    .A(execution_unit_0.inst_ad_0_ ),
    .B(execution_unit_0.inst_type_2_ ),
    .Y(_01367_)
  );
  OAI21X1 _07749_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_alu ),
    .B(_01367_),
    .C(_01366_),
    .Y(_01368_)
  );
  OAI21X1 _07750_ (
    .A(execution_unit_0.inst_type_1_ ),
    .B(_01368_),
    .C(execution_unit_0.alu_0.exec_cycle ),
    .Y(_01369_)
  );
  NAND2X1 _07751_ (
    .A(_01066_),
    .B(_01369_),
    .Y(execution_unit_0.reg_dest_wr )
  );
  OR2X1 _07752_ (
    .A(execution_unit_0.inst_as_1_ ),
    .B(_01278_),
    .Y(_01370_)
  );
  NOR2X1 _07753_ (
    .A(_01152_),
    .B(_01370_),
    .Y(_01371_)
  );
  NOR2X1 _07754_ (
    .A(_01280_),
    .B(_01371_),
    .Y(_01372_)
  );
  OAI21X1 _07755_ (
    .A(execution_unit_0.inst_irq_rst ),
    .B(_01112_),
    .C(_01372_),
    .Y(execution_unit_0.reg_sp_wr )
  );
  OAI21X1 _07756_ (
    .A(_01028_),
    .B(_01069_),
    .C(_01262_),
    .Y(execution_unit_0.reg_pc_call )
  );
  AOI22X1 _07757_ (
    .A(execution_unit_0.inst_as_3_ ),
    .B(exec_done),
    .C(execution_unit_0.alu_0.exec_cycle ),
    .D(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_01373_)
  );
  OAI21X1 _07758_ (
    .A(_01037_),
    .B(_01073_),
    .C(_01373_),
    .Y(execution_unit_0.reg_incr )
  );
  AOI21X1 _07759_ (
    .A(dbg_0.UNUSED_eu_mab_0_ ),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01118_),
    .Y(dbg_0.UNUSED_eu_mb_wr_0_ )
  );
  AOI21X1 _07760_ (
    .A(_01040_),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(_01118_),
    .Y(dbg_0.UNUSED_eu_mb_wr_1_ )
  );
  DFFSR _07761_ (
    .CLK(dco_clk),
    .D(_00991_),
    .Q(execution_unit_0.mdb_in_buf_0_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07762_ (
    .CLK(dco_clk),
    .D(_00998_),
    .Q(execution_unit_0.mdb_in_buf_1_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07763_ (
    .CLK(dco_clk),
    .D(_00999_),
    .Q(execution_unit_0.mdb_in_buf_2_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07764_ (
    .CLK(dco_clk),
    .D(_01000_),
    .Q(execution_unit_0.mdb_in_buf_3_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07765_ (
    .CLK(dco_clk),
    .D(_01001_),
    .Q(execution_unit_0.mdb_in_buf_4_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07766_ (
    .CLK(dco_clk),
    .D(_01002_),
    .Q(execution_unit_0.mdb_in_buf_5_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07767_ (
    .CLK(dco_clk),
    .D(_01003_),
    .Q(execution_unit_0.mdb_in_buf_6_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07768_ (
    .CLK(dco_clk),
    .D(_01004_),
    .Q(execution_unit_0.mdb_in_buf_7_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07769_ (
    .CLK(dco_clk),
    .D(_01005_),
    .Q(execution_unit_0.mdb_in_buf_8_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07770_ (
    .CLK(dco_clk),
    .D(_01006_),
    .Q(execution_unit_0.mdb_in_buf_9_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07771_ (
    .CLK(dco_clk),
    .D(_00992_),
    .Q(execution_unit_0.mdb_in_buf_10_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07772_ (
    .CLK(dco_clk),
    .D(_00993_),
    .Q(execution_unit_0.mdb_in_buf_11_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07773_ (
    .CLK(dco_clk),
    .D(_00994_),
    .Q(execution_unit_0.mdb_in_buf_12_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07774_ (
    .CLK(dco_clk),
    .D(_00995_),
    .Q(execution_unit_0.mdb_in_buf_13_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07775_ (
    .CLK(dco_clk),
    .D(_00996_),
    .Q(execution_unit_0.mdb_in_buf_14_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07776_ (
    .CLK(dco_clk),
    .D(_00997_),
    .Q(execution_unit_0.mdb_in_buf_15_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07777_ (
    .CLK(dco_clk),
    .D(_01008_),
    .Q(execution_unit_0.mdb_in_buf_valid ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07778_ (
    .CLK(dco_clk),
    .D(_01007_),
    .Q(execution_unit_0.mdb_in_buf_en ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07779_ (
    .CLK(dco_clk),
    .D(_00990_),
    .Q(execution_unit_0.mab_lsb ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07780_ (
    .CLK(dco_clk),
    .D(_01009_),
    .Q(eu_mdb_out_0_),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07781_ (
    .CLK(dco_clk),
    .D(_01016_),
    .Q(eu_mdb_out_1_),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07782_ (
    .CLK(dco_clk),
    .D(_01017_),
    .Q(eu_mdb_out_2_),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07783_ (
    .CLK(dco_clk),
    .D(_01018_),
    .Q(eu_mdb_out_3_),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07784_ (
    .CLK(dco_clk),
    .D(_01019_),
    .Q(eu_mdb_out_4_),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07785_ (
    .CLK(dco_clk),
    .D(_01020_),
    .Q(eu_mdb_out_5_),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07786_ (
    .CLK(dco_clk),
    .D(_01021_),
    .Q(eu_mdb_out_6_),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07787_ (
    .CLK(dco_clk),
    .D(_01022_),
    .Q(eu_mdb_out_7_),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07788_ (
    .CLK(dco_clk),
    .D(_01023_),
    .Q(execution_unit_0.mdb_out_nxt_8_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07789_ (
    .CLK(dco_clk),
    .D(_01024_),
    .Q(execution_unit_0.mdb_out_nxt_9_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07790_ (
    .CLK(dco_clk),
    .D(_01010_),
    .Q(execution_unit_0.mdb_out_nxt_10_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07791_ (
    .CLK(dco_clk),
    .D(_01011_),
    .Q(execution_unit_0.mdb_out_nxt_11_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07792_ (
    .CLK(dco_clk),
    .D(_01012_),
    .Q(execution_unit_0.mdb_out_nxt_12_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07793_ (
    .CLK(dco_clk),
    .D(_01013_),
    .Q(execution_unit_0.mdb_out_nxt_13_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07794_ (
    .CLK(dco_clk),
    .D(_01014_),
    .Q(execution_unit_0.mdb_out_nxt_14_ ),
    .R(_01025_),
    .S(1'h1)
  );
  DFFSR _07795_ (
    .CLK(dco_clk),
    .D(_01015_),
    .Q(execution_unit_0.mdb_out_nxt_15_ ),
    .R(_01025_),
    .S(1'h1)
  );
  INVX1 _07796_ (
    .A(execution_unit_0.alu_0.exec_cycle ),
    .Y(_01919_)
  );
  INVX1 _07797_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .Y(_01374_)
  );
  INVX1 _07798_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01375_)
  );
  INVX1 _07799_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01376_)
  );
  INVX1 _07800_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01377_)
  );
  INVX1 _07801_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .Y(_01378_)
  );
  INVX1 _07802_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01379_)
  );
  INVX1 _07803_ (
    .A(execution_unit_0.alu_0.inst_jmp_4_ ),
    .Y(_01380_)
  );
  INVX1 _07804_ (
    .A(execution_unit_0.alu_0.inst_jmp_1_ ),
    .Y(_01381_)
  );
  INVX1 _07805_ (
    .A(execution_unit_0.alu_0.alu_shift_3_ ),
    .Y(_01382_)
  );
  INVX1 _07806_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .Y(_01383_)
  );
  INVX1 _07807_ (
    .A(execution_unit_0.alu_0.op_dst_15_ ),
    .Y(_01384_)
  );
  OR2X1 _07808_ (
    .A(cpu_halt_st),
    .B(execution_unit_0.alu_0.inst_so_7_ ),
    .Y(_01385_)
  );
  NOR2X1 _07809_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01385_),
    .Y(_01386_)
  );
  OR2X1 _07810_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01385_),
    .Y(_01387_)
  );
  AND2X1 _07811_ (
    .A(execution_unit_0.alu_0.inst_alu_0_ ),
    .B(execution_unit_0.alu_0.exec_cycle ),
    .Y(_01388_)
  );
  NAND2X1 _07812_ (
    .A(execution_unit_0.alu_0.inst_alu_0_ ),
    .B(execution_unit_0.alu_0.exec_cycle ),
    .Y(_01389_)
  );
  XNOR2X1 _07813_ (
    .A(execution_unit_0.alu_0.alu_swpb_8_ ),
    .B(_01389_),
    .Y(_01390_)
  );
  AND2X1 _07814_ (
    .A(execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01390_),
    .Y(_01391_)
  );
  NAND2X1 _07815_ (
    .A(execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01390_),
    .Y(_01392_)
  );
  NAND2X1 _07816_ (
    .A(execution_unit_0.alu_0.status_1_ ),
    .B(execution_unit_0.alu_0.inst_jmp_0_ ),
    .Y(_01393_)
  );
  OAI21X1 _07817_ (
    .A(_01381_),
    .B(execution_unit_0.alu_0.status_1_ ),
    .C(_01393_),
    .Y(_01394_)
  );
  MUX2X1 _07818_ (
    .A(execution_unit_0.alu_0.inst_jmp_2_ ),
    .B(execution_unit_0.alu_0.inst_jmp_3_ ),
    .S(execution_unit_0.alu_0.status_0_ ),
    .Y(_01395_)
  );
  OAI21X1 _07819_ (
    .A(execution_unit_0.alu_0.status_2_ ),
    .B(_01380_),
    .C(_01395_),
    .Y(_01396_)
  );
  NOR2X1 _07820_ (
    .A(_01394_),
    .B(_01396_),
    .Y(_01397_)
  );
  XOR2X1 _07821_ (
    .A(execution_unit_0.alu_0.status_3_ ),
    .B(execution_unit_0.alu_0.status_2_ ),
    .Y(_01398_)
  );
  MUX2X1 _07822_ (
    .A(execution_unit_0.alu_0.inst_jmp_5_ ),
    .B(execution_unit_0.alu_0.inst_jmp_6_ ),
    .S(_01398_),
    .Y(_01399_)
  );
  AND2X1 _07823_ (
    .A(_01397_),
    .B(_01399_),
    .Y(_01400_)
  );
  NAND2X1 _07824_ (
    .A(_01397_),
    .B(_01399_),
    .Y(_01401_)
  );
  AOI21X1 _07825_ (
    .A(_01390_),
    .B(_01400_),
    .C(execution_unit_0.alu_0.op_dst_0_ ),
    .Y(_01402_)
  );
  AOI21X1 _07826_ (
    .A(_01391_),
    .B(_01400_),
    .C(_01402_),
    .Y(dbg_0.UNUSED_eu_mab_0_ )
  );
  AOI21X1 _07827_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(execution_unit_0.alu_0.inst_alu_2_ ),
    .C(execution_unit_0.alu_0.inst_alu_1_ ),
    .Y(_01403_)
  );
  NOR2X1 _07828_ (
    .A(_01919_),
    .B(_01403_),
    .Y(_01404_)
  );
  NAND2X1 _07829_ (
    .A(dbg_0.UNUSED_eu_mab_0_ ),
    .B(_01404_),
    .Y(_01405_)
  );
  OR2X1 _07830_ (
    .A(dbg_0.UNUSED_eu_mab_0_ ),
    .B(_01404_),
    .Y(_01406_)
  );
  NOR2X1 _07831_ (
    .A(execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01390_),
    .Y(_01407_)
  );
  OR2X1 _07832_ (
    .A(execution_unit_0.alu_0.op_dst_0_ ),
    .B(_01390_),
    .Y(_01408_)
  );
  NAND2X1 _07833_ (
    .A(_01392_),
    .B(_01408_),
    .Y(_01409_)
  );
  XNOR2X1 _07834_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(_01409_),
    .Y(_01410_)
  );
  NOR2X1 _07835_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(execution_unit_0.alu_0.inst_so_3_ ),
    .Y(_01411_)
  );
  NOR2X1 _07836_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01412_)
  );
  NAND2X1 _07837_ (
    .A(_01377_),
    .B(_01412_),
    .Y(_01413_)
  );
  NAND2X1 _07838_ (
    .A(_01374_),
    .B(_01411_),
    .Y(_01414_)
  );
  NOR2X1 _07839_ (
    .A(_01413_),
    .B(_01414_),
    .Y(_01415_)
  );
  AOI21X1 _07840_ (
    .A(execution_unit_0.alu_0.alu_shift_0_ ),
    .B(execution_unit_0.alu_0.inst_alu_10_ ),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01416_)
  );
  AOI22X1 _07841_ (
    .A(execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(execution_unit_0.alu_0.inst_so_1_ ),
    .C(execution_unit_0.alu_0.inst_so_3_ ),
    .D(execution_unit_0.alu_0.alu_swpb_8_ ),
    .Y(_01417_)
  );
  NAND2X1 _07842_ (
    .A(_01416_),
    .B(_01417_),
    .Y(_01418_)
  );
  AOI21X1 _07843_ (
    .A(_01390_),
    .B(_01415_),
    .C(_01418_),
    .Y(_01419_)
  );
  OAI21X1 _07844_ (
    .A(_01376_),
    .B(_01392_),
    .C(_01419_),
    .Y(_01420_)
  );
  AOI21X1 _07845_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01408_),
    .C(_01420_),
    .Y(_01421_)
  );
  OAI21X1 _07846_ (
    .A(_01374_),
    .B(_01409_),
    .C(_01421_),
    .Y(_01422_)
  );
  OAI21X1 _07847_ (
    .A(_01379_),
    .B(_01410_),
    .C(_01422_),
    .Y(_01423_)
  );
  NAND3X1 _07848_ (
    .A(_01387_),
    .B(_01405_),
    .C(_01406_),
    .Y(_01424_)
  );
  OAI21X1 _07849_ (
    .A(_01387_),
    .B(_01423_),
    .C(_01424_),
    .Y(execution_unit_0.alu_0.alu_out_0_ )
  );
  XNOR2X1 _07850_ (
    .A(execution_unit_0.alu_0.alu_shift_0_ ),
    .B(_01389_),
    .Y(_01425_)
  );
  AND2X1 _07851_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01425_),
    .Y(_01426_)
  );
  NAND2X1 _07852_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01425_),
    .Y(_01427_)
  );
  NOR2X1 _07853_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01425_),
    .Y(_01428_)
  );
  NOR2X1 _07854_ (
    .A(_01426_),
    .B(_01428_),
    .Y(_01429_)
  );
  OR2X1 _07855_ (
    .A(_01426_),
    .B(_01428_),
    .Y(_01430_)
  );
  NAND3X1 _07856_ (
    .A(_01391_),
    .B(_01400_),
    .C(_01429_),
    .Y(_01431_)
  );
  NAND3X1 _07857_ (
    .A(_01392_),
    .B(_01400_),
    .C(_01430_),
    .Y(_01432_)
  );
  AND2X1 _07858_ (
    .A(_01431_),
    .B(_01432_),
    .Y(_01433_)
  );
  OAI21X1 _07859_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01400_),
    .C(_01433_),
    .Y(_01434_)
  );
  INVX1 _07860_ (
    .A(_01434_),
    .Y(dbg_0.UNUSED_eu_mab_1_ )
  );
  OR2X1 _07861_ (
    .A(_01405_),
    .B(_01434_),
    .Y(_01435_)
  );
  OAI21X1 _07862_ (
    .A(_01405_),
    .B(_01434_),
    .C(_01387_),
    .Y(_01436_)
  );
  AOI21X1 _07863_ (
    .A(_01405_),
    .B(_01434_),
    .C(_01436_),
    .Y(_01437_)
  );
  AOI21X1 _07864_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(_01408_),
    .C(_01391_),
    .Y(_01438_)
  );
  OAI21X1 _07865_ (
    .A(_01378_),
    .B(_01407_),
    .C(_01392_),
    .Y(_01439_)
  );
  XNOR2X1 _07866_ (
    .A(_01430_),
    .B(_01438_),
    .Y(_01440_)
  );
  INVX1 _07867_ (
    .A(_01440_),
    .Y(_01441_)
  );
  AOI21X1 _07868_ (
    .A(_01429_),
    .B(_01439_),
    .C(_01426_),
    .Y(_01442_)
  );
  OAI21X1 _07869_ (
    .A(_01430_),
    .B(_01438_),
    .C(_01427_),
    .Y(_01443_)
  );
  XNOR2X1 _07870_ (
    .A(execution_unit_0.alu_0.alu_shift_1_ ),
    .B(_01389_),
    .Y(_01444_)
  );
  AND2X1 _07871_ (
    .A(execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01444_),
    .Y(_01445_)
  );
  NAND2X1 _07872_ (
    .A(execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01444_),
    .Y(_01446_)
  );
  OR2X1 _07873_ (
    .A(execution_unit_0.alu_0.op_dst_2_ ),
    .B(_01444_),
    .Y(_01447_)
  );
  INVX1 _07874_ (
    .A(_01447_),
    .Y(_01448_)
  );
  NAND2X1 _07875_ (
    .A(_01446_),
    .B(_01447_),
    .Y(_01449_)
  );
  XNOR2X1 _07876_ (
    .A(_01443_),
    .B(_01449_),
    .Y(_01450_)
  );
  NOR2X1 _07877_ (
    .A(_01441_),
    .B(_01450_),
    .Y(_01451_)
  );
  OR2X1 _07878_ (
    .A(_01441_),
    .B(_01450_),
    .Y(_01452_)
  );
  AOI21X1 _07879_ (
    .A(_01443_),
    .B(_01447_),
    .C(_01445_),
    .Y(_01453_)
  );
  OAI21X1 _07880_ (
    .A(_01442_),
    .B(_01448_),
    .C(_01446_),
    .Y(_01454_)
  );
  XNOR2X1 _07881_ (
    .A(execution_unit_0.alu_0.alu_shift_2_ ),
    .B(_01389_),
    .Y(_01455_)
  );
  AND2X1 _07882_ (
    .A(execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01455_),
    .Y(_01456_)
  );
  NAND2X1 _07883_ (
    .A(execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01455_),
    .Y(_01457_)
  );
  OR2X1 _07884_ (
    .A(execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01455_),
    .Y(_01458_)
  );
  INVX1 _07885_ (
    .A(_01458_),
    .Y(_01459_)
  );
  NAND2X1 _07886_ (
    .A(_01457_),
    .B(_01458_),
    .Y(_01460_)
  );
  XNOR2X1 _07887_ (
    .A(_01454_),
    .B(_01460_),
    .Y(_01461_)
  );
  XNOR2X1 _07888_ (
    .A(_01453_),
    .B(_01460_),
    .Y(_01462_)
  );
  OAI21X1 _07889_ (
    .A(_01454_),
    .B(_01456_),
    .C(_01458_),
    .Y(_01463_)
  );
  AOI21X1 _07890_ (
    .A(_01453_),
    .B(_01457_),
    .C(_01459_),
    .Y(_01464_)
  );
  AOI21X1 _07891_ (
    .A(_01452_),
    .B(_01461_),
    .C(_01464_),
    .Y(_01465_)
  );
  OAI21X1 _07892_ (
    .A(_01451_),
    .B(_01462_),
    .C(_01463_),
    .Y(_01466_)
  );
  NAND2X1 _07893_ (
    .A(_01440_),
    .B(_01466_),
    .Y(_01467_)
  );
  AOI21X1 _07894_ (
    .A(_01441_),
    .B(_01465_),
    .C(_01379_),
    .Y(_01468_)
  );
  OAI21X1 _07895_ (
    .A(execution_unit_0.alu_0.op_dst_1_ ),
    .B(_01425_),
    .C(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01469_)
  );
  NAND2X1 _07896_ (
    .A(_01415_),
    .B(_01425_),
    .Y(_01470_)
  );
  AOI22X1 _07897_ (
    .A(execution_unit_0.alu_0.alu_shift_0_ ),
    .B(execution_unit_0.alu_0.inst_so_3_ ),
    .C(_01426_),
    .D(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01471_)
  );
  OAI21X1 _07898_ (
    .A(_01374_),
    .B(_01430_),
    .C(_01471_),
    .Y(_01472_)
  );
  AOI22X1 _07899_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_8_ ),
    .C(execution_unit_0.alu_0.alu_shift_1_ ),
    .D(execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01473_)
  );
  NAND3X1 _07900_ (
    .A(_01469_),
    .B(_01470_),
    .C(_01473_),
    .Y(_01474_)
  );
  OR2X1 _07901_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01474_),
    .Y(_01475_)
  );
  OAI21X1 _07902_ (
    .A(_01472_),
    .B(_01475_),
    .C(_01386_),
    .Y(_01476_)
  );
  AOI21X1 _07903_ (
    .A(_01467_),
    .B(_01468_),
    .C(_01476_),
    .Y(_01477_)
  );
  NOR2X1 _07904_ (
    .A(_01437_),
    .B(_01477_),
    .Y(_01478_)
  );
  INVX1 _07905_ (
    .A(_01478_),
    .Y(execution_unit_0.alu_0.alu_out_1_ )
  );
  OAI21X1 _07906_ (
    .A(_01401_),
    .B(_01427_),
    .C(_01431_),
    .Y(_01479_)
  );
  AOI21X1 _07907_ (
    .A(_01400_),
    .B(_01444_),
    .C(execution_unit_0.alu_0.op_dst_2_ ),
    .Y(_01480_)
  );
  AOI21X1 _07908_ (
    .A(_01400_),
    .B(_01445_),
    .C(_01480_),
    .Y(_01481_)
  );
  XNOR2X1 _07909_ (
    .A(_01479_),
    .B(_01481_),
    .Y(_01482_)
  );
  INVX1 _07910_ (
    .A(_01482_),
    .Y(dbg_0.UNUSED_eu_mab_2_ )
  );
  AND2X1 _07911_ (
    .A(_01435_),
    .B(_01482_),
    .Y(_01483_)
  );
  NOR2X1 _07912_ (
    .A(_01435_),
    .B(_01482_),
    .Y(_01484_)
  );
  OAI21X1 _07913_ (
    .A(_01435_),
    .B(_01482_),
    .C(_01387_),
    .Y(_01485_)
  );
  OAI21X1 _07914_ (
    .A(_01452_),
    .B(_01463_),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01486_)
  );
  AOI21X1 _07915_ (
    .A(_01450_),
    .B(_01467_),
    .C(_01486_),
    .Y(_01487_)
  );
  AOI22X1 _07916_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_1_ ),
    .C(execution_unit_0.alu_0.alu_shift_2_ ),
    .D(execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01488_)
  );
  OAI21X1 _07917_ (
    .A(_01376_),
    .B(_01446_),
    .C(_01488_),
    .Y(_01489_)
  );
  AOI21X1 _07918_ (
    .A(_01415_),
    .B(_01444_),
    .C(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01490_)
  );
  NOR2X1 _07919_ (
    .A(_01448_),
    .B(_01490_),
    .Y(_01491_)
  );
  OR2X1 _07920_ (
    .A(_01489_),
    .B(_01491_),
    .Y(_01492_)
  );
  AOI21X1 _07921_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_9_ ),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01493_)
  );
  OAI21X1 _07922_ (
    .A(_01374_),
    .B(_01449_),
    .C(_01493_),
    .Y(_01494_)
  );
  OAI21X1 _07923_ (
    .A(_01492_),
    .B(_01494_),
    .C(_01386_),
    .Y(_01495_)
  );
  OAI22X1 _07924_ (
    .A(_01483_),
    .B(_01485_),
    .C(_01487_),
    .D(_01495_),
    .Y(execution_unit_0.alu_0.alu_out_2_ )
  );
  AOI22X1 _07925_ (
    .A(_01400_),
    .B(_01445_),
    .C(_01479_),
    .D(_01481_),
    .Y(_01496_)
  );
  OAI21X1 _07926_ (
    .A(execution_unit_0.alu_0.op_dst_3_ ),
    .B(_01400_),
    .C(_01458_),
    .Y(_01497_)
  );
  AOI21X1 _07927_ (
    .A(_01400_),
    .B(_01456_),
    .C(_01497_),
    .Y(_01498_)
  );
  XNOR2X1 _07928_ (
    .A(_01496_),
    .B(_01498_),
    .Y(dbg_0.UNUSED_eu_mab_3_ )
  );
  NAND2X1 _07929_ (
    .A(_01484_),
    .B(dbg_0.UNUSED_eu_mab_3_ ),
    .Y(_01499_)
  );
  XNOR2X1 _07930_ (
    .A(_01484_),
    .B(dbg_0.UNUSED_eu_mab_3_ ),
    .Y(_01500_)
  );
  OAI21X1 _07931_ (
    .A(_01451_),
    .B(_01463_),
    .C(_01462_),
    .Y(_01501_)
  );
  AND2X1 _07932_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01501_),
    .Y(_01502_)
  );
  OAI21X1 _07933_ (
    .A(_01451_),
    .B(_01462_),
    .C(_01502_),
    .Y(_01503_)
  );
  NAND2X1 _07934_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01386_),
    .Y(_01504_)
  );
  AOI22X1 _07935_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_2_ ),
    .C(execution_unit_0.alu_0.alu_shift_10_ ),
    .D(execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01505_)
  );
  OAI21X1 _07936_ (
    .A(_01377_),
    .B(_01382_),
    .C(_01505_),
    .Y(_01506_)
  );
  AOI22X1 _07937_ (
    .A(_01415_),
    .B(_01455_),
    .C(_01458_),
    .D(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01507_)
  );
  AOI21X1 _07938_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01456_),
    .C(_01506_),
    .Y(_01508_)
  );
  NAND2X1 _07939_ (
    .A(_01507_),
    .B(_01508_),
    .Y(_01509_)
  );
  OAI21X1 _07940_ (
    .A(_01374_),
    .B(_01460_),
    .C(_01386_),
    .Y(_01510_)
  );
  OAI21X1 _07941_ (
    .A(_01509_),
    .B(_01510_),
    .C(_01504_),
    .Y(_01511_)
  );
  AOI22X1 _07942_ (
    .A(_01387_),
    .B(_01500_),
    .C(_01503_),
    .D(_01511_),
    .Y(execution_unit_0.alu_0.alu_out_3_ )
  );
  XNOR2X1 _07943_ (
    .A(_01382_),
    .B(_01388_),
    .Y(_01512_)
  );
  AND2X1 _07944_ (
    .A(execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01512_),
    .Y(_01513_)
  );
  NAND2X1 _07945_ (
    .A(execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01512_),
    .Y(_01514_)
  );
  NAND2X1 _07946_ (
    .A(_01400_),
    .B(_01512_),
    .Y(_01515_)
  );
  XOR2X1 _07947_ (
    .A(execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01515_),
    .Y(_01516_)
  );
  INVX1 _07948_ (
    .A(_01516_),
    .Y(_01517_)
  );
  OAI22X1 _07949_ (
    .A(_01401_),
    .B(_01457_),
    .C(_01496_),
    .D(_01497_),
    .Y(_01518_)
  );
  XNOR2X1 _07950_ (
    .A(_01517_),
    .B(_01518_),
    .Y(_01519_)
  );
  INVX1 _07951_ (
    .A(_01519_),
    .Y(dbg_0.UNUSED_eu_mab_4_ )
  );
  AND2X1 _07952_ (
    .A(_01499_),
    .B(_01519_),
    .Y(_01520_)
  );
  NOR2X1 _07953_ (
    .A(_01499_),
    .B(_01519_),
    .Y(_01521_)
  );
  NOR2X1 _07954_ (
    .A(execution_unit_0.alu_0.op_dst_4_ ),
    .B(_01512_),
    .Y(_01522_)
  );
  NOR2X1 _07955_ (
    .A(_01513_),
    .B(_01522_),
    .Y(_01523_)
  );
  OR2X1 _07956_ (
    .A(_01513_),
    .B(_01522_),
    .Y(_01524_)
  );
  NOR3X1 _07957_ (
    .A(_01451_),
    .B(_01462_),
    .C(_01463_),
    .Y(_01525_)
  );
  NAND3X1 _07958_ (
    .A(_01452_),
    .B(_01461_),
    .C(_01464_),
    .Y(_01526_)
  );
  NOR3X1 _07959_ (
    .A(_01465_),
    .B(_01524_),
    .C(_01525_),
    .Y(_01527_)
  );
  NAND3X1 _07960_ (
    .A(_01466_),
    .B(_01523_),
    .C(_01526_),
    .Y(_01528_)
  );
  AOI21X1 _07961_ (
    .A(_01466_),
    .B(_01526_),
    .C(_01523_),
    .Y(_01529_)
  );
  OAI21X1 _07962_ (
    .A(_01527_),
    .B(_01529_),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01530_)
  );
  NOR2X1 _07963_ (
    .A(_01375_),
    .B(_01522_),
    .Y(_01531_)
  );
  AOI21X1 _07964_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_4_ ),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01532_)
  );
  AOI22X1 _07965_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_3_ ),
    .C(execution_unit_0.alu_0.alu_shift_11_ ),
    .D(execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01533_)
  );
  NAND2X1 _07966_ (
    .A(_01532_),
    .B(_01533_),
    .Y(_01534_)
  );
  AOI21X1 _07967_ (
    .A(_01415_),
    .B(_01512_),
    .C(_01534_),
    .Y(_01535_)
  );
  OAI21X1 _07968_ (
    .A(_01376_),
    .B(_01514_),
    .C(_01535_),
    .Y(_01536_)
  );
  NOR2X1 _07969_ (
    .A(_01531_),
    .B(_01536_),
    .Y(_01537_)
  );
  OAI21X1 _07970_ (
    .A(_01374_),
    .B(_01524_),
    .C(_01537_),
    .Y(_01538_)
  );
  OAI21X1 _07971_ (
    .A(_01499_),
    .B(_01519_),
    .C(_01387_),
    .Y(_01539_)
  );
  NAND3X1 _07972_ (
    .A(_01386_),
    .B(_01530_),
    .C(_01538_),
    .Y(_01540_)
  );
  OAI21X1 _07973_ (
    .A(_01520_),
    .B(_01539_),
    .C(_01540_),
    .Y(execution_unit_0.alu_0.alu_out_4_ )
  );
  AOI22X1 _07974_ (
    .A(_01400_),
    .B(_01513_),
    .C(_01517_),
    .D(_01518_),
    .Y(_01541_)
  );
  XNOR2X1 _07975_ (
    .A(execution_unit_0.alu_0.alu_shift_4_ ),
    .B(_01389_),
    .Y(_01542_)
  );
  AND2X1 _07976_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01542_),
    .Y(_01543_)
  );
  NAND2X1 _07977_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01542_),
    .Y(_01544_)
  );
  NAND2X1 _07978_ (
    .A(_01400_),
    .B(_01542_),
    .Y(_01545_)
  );
  XOR2X1 _07979_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01545_),
    .Y(_01546_)
  );
  XOR2X1 _07980_ (
    .A(_01541_),
    .B(_01546_),
    .Y(dbg_0.UNUSED_eu_mab_5_ )
  );
  NOR2X1 _07981_ (
    .A(_01521_),
    .B(dbg_0.UNUSED_eu_mab_5_ ),
    .Y(_01547_)
  );
  NAND2X1 _07982_ (
    .A(_01521_),
    .B(dbg_0.UNUSED_eu_mab_5_ ),
    .Y(_01548_)
  );
  OAI21X1 _07983_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01385_),
    .C(_01548_),
    .Y(_01549_)
  );
  XNOR2X1 _07984_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01542_),
    .Y(_01550_)
  );
  INVX1 _07985_ (
    .A(_01550_),
    .Y(_01551_)
  );
  AOI21X1 _07986_ (
    .A(_01514_),
    .B(_01528_),
    .C(_01550_),
    .Y(_01552_)
  );
  OAI21X1 _07987_ (
    .A(_01513_),
    .B(_01527_),
    .C(_01551_),
    .Y(_01553_)
  );
  NAND3X1 _07988_ (
    .A(_01514_),
    .B(_01528_),
    .C(_01550_),
    .Y(_01554_)
  );
  AND2X1 _07989_ (
    .A(_01553_),
    .B(_01554_),
    .Y(_01555_)
  );
  XNOR2X1 _07990_ (
    .A(execution_unit_0.alu_0.alu_shift_5_ ),
    .B(_01389_),
    .Y(_01556_)
  );
  AND2X1 _07991_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01556_),
    .Y(_01557_)
  );
  NAND2X1 _07992_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01556_),
    .Y(_01558_)
  );
  XNOR2X1 _07993_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01556_),
    .Y(_01559_)
  );
  INVX1 _07994_ (
    .A(_01559_),
    .Y(_01560_)
  );
  AOI21X1 _07995_ (
    .A(_01544_),
    .B(_01553_),
    .C(_01559_),
    .Y(_01561_)
  );
  OAI21X1 _07996_ (
    .A(_01543_),
    .B(_01552_),
    .C(_01560_),
    .Y(_01562_)
  );
  NAND3X1 _07997_ (
    .A(_01544_),
    .B(_01553_),
    .C(_01559_),
    .Y(_01563_)
  );
  NAND2X1 _07998_ (
    .A(_01562_),
    .B(_01563_),
    .Y(_01564_)
  );
  AOI21X1 _07999_ (
    .A(_01562_),
    .B(_01563_),
    .C(_01555_),
    .Y(_01565_)
  );
  XNOR2X1 _08000_ (
    .A(execution_unit_0.alu_0.alu_shift_6_ ),
    .B(_01389_),
    .Y(_01566_)
  );
  AND2X1 _08001_ (
    .A(execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01566_),
    .Y(_01567_)
  );
  NOR2X1 _08002_ (
    .A(execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01566_),
    .Y(_01568_)
  );
  NOR2X1 _08003_ (
    .A(_01567_),
    .B(_01568_),
    .Y(_01569_)
  );
  INVX1 _08004_ (
    .A(_01569_),
    .Y(_01570_)
  );
  NAND3X1 _08005_ (
    .A(_01558_),
    .B(_01562_),
    .C(_01569_),
    .Y(_01571_)
  );
  OAI21X1 _08006_ (
    .A(_01557_),
    .B(_01561_),
    .C(_01570_),
    .Y(_01572_)
  );
  NAND2X1 _08007_ (
    .A(_01571_),
    .B(_01572_),
    .Y(_01573_)
  );
  AOI21X1 _08008_ (
    .A(_01571_),
    .B(_01572_),
    .C(_01565_),
    .Y(_01574_)
  );
  INVX1 _08009_ (
    .A(_01574_),
    .Y(_01575_)
  );
  AOI21X1 _08010_ (
    .A(_01558_),
    .B(_01562_),
    .C(_01568_),
    .Y(_01576_)
  );
  NOR2X1 _08011_ (
    .A(_01567_),
    .B(_01576_),
    .Y(_01577_)
  );
  NAND2X1 _08012_ (
    .A(_01575_),
    .B(_01577_),
    .Y(_01578_)
  );
  AOI21X1 _08013_ (
    .A(_01575_),
    .B(_01577_),
    .C(_01555_),
    .Y(_01579_)
  );
  XNOR2X1 _08014_ (
    .A(_01555_),
    .B(_01578_),
    .Y(_01580_)
  );
  NOR2X1 _08015_ (
    .A(_01374_),
    .B(_01550_),
    .Y(_01581_)
  );
  OAI21X1 _08016_ (
    .A(execution_unit_0.alu_0.op_dst_5_ ),
    .B(_01542_),
    .C(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01582_)
  );
  NAND2X1 _08017_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01543_),
    .Y(_01583_)
  );
  AOI21X1 _08018_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_5_ ),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01584_)
  );
  AOI22X1 _08019_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_4_ ),
    .C(execution_unit_0.alu_0.alu_shift_12_ ),
    .D(execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01585_)
  );
  NAND2X1 _08020_ (
    .A(_01584_),
    .B(_01585_),
    .Y(_01586_)
  );
  AOI21X1 _08021_ (
    .A(_01415_),
    .B(_01542_),
    .C(_01586_),
    .Y(_01587_)
  );
  NAND3X1 _08022_ (
    .A(_01582_),
    .B(_01583_),
    .C(_01587_),
    .Y(_01588_)
  );
  OAI21X1 _08023_ (
    .A(_01581_),
    .B(_01588_),
    .C(_01386_),
    .Y(_01589_)
  );
  AOI21X1 _08024_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01580_),
    .C(_01589_),
    .Y(_01590_)
  );
  INVX1 _08025_ (
    .A(_01590_),
    .Y(_01591_)
  );
  OAI21X1 _08026_ (
    .A(_01547_),
    .B(_01549_),
    .C(_01591_),
    .Y(execution_unit_0.alu_0.alu_out_5_ )
  );
  OAI22X1 _08027_ (
    .A(_01401_),
    .B(_01544_),
    .C(_01546_),
    .D(_01541_),
    .Y(_01592_)
  );
  NAND2X1 _08028_ (
    .A(_01400_),
    .B(_01556_),
    .Y(_01593_)
  );
  XOR2X1 _08029_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01593_),
    .Y(_01594_)
  );
  INVX1 _08030_ (
    .A(_01594_),
    .Y(_01595_)
  );
  NAND2X1 _08031_ (
    .A(_01592_),
    .B(_01595_),
    .Y(_01596_)
  );
  XNOR2X1 _08032_ (
    .A(_01592_),
    .B(_01595_),
    .Y(_01597_)
  );
  INVX1 _08033_ (
    .A(_01597_),
    .Y(dbg_0.UNUSED_eu_mab_6_ )
  );
  NOR2X1 _08034_ (
    .A(_01548_),
    .B(_01597_),
    .Y(_01598_)
  );
  XNOR2X1 _08035_ (
    .A(_01548_),
    .B(_01597_),
    .Y(_01599_)
  );
  NOR2X1 _08036_ (
    .A(_01374_),
    .B(_01559_),
    .Y(_01600_)
  );
  OAI21X1 _08037_ (
    .A(execution_unit_0.alu_0.op_dst_6_ ),
    .B(_01556_),
    .C(execution_unit_0.alu_0.inst_alu_5_ ),
    .Y(_01601_)
  );
  AOI22X1 _08038_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_5_ ),
    .C(execution_unit_0.alu_0.alu_shift_13_ ),
    .D(execution_unit_0.alu_0.inst_so_1_ ),
    .Y(_01602_)
  );
  NAND2X1 _08039_ (
    .A(_01386_),
    .B(_01602_),
    .Y(_01603_)
  );
  AOI21X1 _08040_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_6_ ),
    .C(_01603_),
    .Y(_01604_)
  );
  AOI22X1 _08041_ (
    .A(_01415_),
    .B(_01556_),
    .C(_01557_),
    .D(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01605_)
  );
  NAND3X1 _08042_ (
    .A(_01601_),
    .B(_01604_),
    .C(_01605_),
    .Y(_01606_)
  );
  OAI21X1 _08043_ (
    .A(_01600_),
    .B(_01606_),
    .C(_01504_),
    .Y(_01607_)
  );
  XNOR2X1 _08044_ (
    .A(_01564_),
    .B(_01579_),
    .Y(_01608_)
  );
  NAND2X1 _08045_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01608_),
    .Y(_01609_)
  );
  AOI22X1 _08046_ (
    .A(_01387_),
    .B(_01599_),
    .C(_01607_),
    .D(_01609_),
    .Y(execution_unit_0.alu_0.alu_out_6_ )
  );
  AOI21X1 _08047_ (
    .A(_01400_),
    .B(_01566_),
    .C(execution_unit_0.alu_0.op_dst_7_ ),
    .Y(_01610_)
  );
  AOI21X1 _08048_ (
    .A(_01400_),
    .B(_01567_),
    .C(_01610_),
    .Y(_01611_)
  );
  OAI21X1 _08049_ (
    .A(_01401_),
    .B(_01558_),
    .C(_01596_),
    .Y(_01612_)
  );
  XOR2X1 _08050_ (
    .A(_01611_),
    .B(_01612_),
    .Y(dbg_0.UNUSED_eu_mab_7_ )
  );
  NAND2X1 _08051_ (
    .A(_01598_),
    .B(dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_01613_)
  );
  XNOR2X1 _08052_ (
    .A(_01598_),
    .B(dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_01614_)
  );
  MUX2X1 _08053_ (
    .A(execution_unit_0.alu_0.alu_shift_6_ ),
    .B(execution_unit_0.alu_0.alu_shift_14_ ),
    .S(execution_unit_0.alu_0.inst_bw ),
    .Y(_01615_)
  );
  NAND2X1 _08054_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(execution_unit_0.alu_0.inst_so_0_ ),
    .Y(_01616_)
  );
  OAI21X1 _08055_ (
    .A(execution_unit_0.alu_0.inst_so_0_ ),
    .B(_01615_),
    .C(_01616_),
    .Y(_01617_)
  );
  NOR2X1 _08056_ (
    .A(_01383_),
    .B(_01617_),
    .Y(_01618_)
  );
  OAI21X1 _08057_ (
    .A(execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(execution_unit_0.alu_0.inst_bw ),
    .C(execution_unit_0.alu_0.inst_alu_10_ ),
    .Y(_01619_)
  );
  NOR2X1 _08058_ (
    .A(_01618_),
    .B(_01619_),
    .Y(_01620_)
  );
  AND2X1 _08059_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(execution_unit_0.alu_0.alu_shift_6_ ),
    .Y(_01621_)
  );
  AOI21X1 _08060_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_14_ ),
    .C(_01621_),
    .Y(_01622_)
  );
  AND2X1 _08061_ (
    .A(_01386_),
    .B(_01622_),
    .Y(_01623_)
  );
  AOI22X1 _08062_ (
    .A(_01415_),
    .B(_01566_),
    .C(_01567_),
    .D(execution_unit_0.alu_0.inst_alu_4_ ),
    .Y(_01624_)
  );
  OAI21X1 _08063_ (
    .A(_01375_),
    .B(_01568_),
    .C(_01623_),
    .Y(_01625_)
  );
  AOI21X1 _08064_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01569_),
    .C(_01625_),
    .Y(_01626_)
  );
  NAND2X1 _08065_ (
    .A(_01624_),
    .B(_01626_),
    .Y(_01627_)
  );
  OAI21X1 _08066_ (
    .A(_01620_),
    .B(_01627_),
    .C(_01504_),
    .Y(_01628_)
  );
  NOR2X1 _08067_ (
    .A(_01565_),
    .B(_01568_),
    .Y(_01629_)
  );
  NOR2X1 _08068_ (
    .A(_01379_),
    .B(_01574_),
    .Y(_01630_)
  );
  OAI21X1 _08069_ (
    .A(_01573_),
    .B(_01629_),
    .C(_01630_),
    .Y(_01631_)
  );
  AOI22X1 _08070_ (
    .A(_01387_),
    .B(_01614_),
    .C(_01628_),
    .D(_01631_),
    .Y(execution_unit_0.alu_0.alu_out_7_ )
  );
  OAI21X1 _08071_ (
    .A(_01557_),
    .B(_01567_),
    .C(_01400_),
    .Y(_01632_)
  );
  OAI22X1 _08072_ (
    .A(_01596_),
    .B(_01610_),
    .C(_01632_),
    .D(_01568_),
    .Y(_01633_)
  );
  NOR2X1 _08073_ (
    .A(_01919_),
    .B(_01383_),
    .Y(_01634_)
  );
  NAND2X1 _08074_ (
    .A(execution_unit_0.alu_0.exec_cycle ),
    .B(execution_unit_0.alu_0.inst_bw ),
    .Y(_01635_)
  );
  OAI21X1 _08075_ (
    .A(execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(_01388_),
    .C(_01635_),
    .Y(_01636_)
  );
  AOI21X1 _08076_ (
    .A(execution_unit_0.alu_0.alu_swpb_0_ ),
    .B(_01388_),
    .C(_01636_),
    .Y(_01637_)
  );
  AND2X1 _08077_ (
    .A(execution_unit_0.alu_0.op_dst_8_ ),
    .B(_01637_),
    .Y(_01638_)
  );
  INVX1 _08078_ (
    .A(_01638_),
    .Y(_01639_)
  );
  NAND2X1 _08079_ (
    .A(_01400_),
    .B(_01638_),
    .Y(_01640_)
  );
  AOI22X1 _08080_ (
    .A(execution_unit_0.alu_0.op_dst_8_ ),
    .B(_01635_),
    .C(_01637_),
    .D(_01400_),
    .Y(_01641_)
  );
  AOI21X1 _08081_ (
    .A(_01400_),
    .B(_01638_),
    .C(_01641_),
    .Y(_01642_)
  );
  NAND2X1 _08082_ (
    .A(_01633_),
    .B(_01642_),
    .Y(_01643_)
  );
  XNOR2X1 _08083_ (
    .A(_01633_),
    .B(_01642_),
    .Y(_01644_)
  );
  INVX1 _08084_ (
    .A(_01644_),
    .Y(dbg_0.UNUSED_eu_mab_8_ )
  );
  AOI21X1 _08085_ (
    .A(execution_unit_0.alu_0.op_dst_8_ ),
    .B(_01635_),
    .C(_01637_),
    .Y(_01645_)
  );
  NOR2X1 _08086_ (
    .A(_01638_),
    .B(_01645_),
    .Y(_01646_)
  );
  XNOR2X1 _08087_ (
    .A(_01574_),
    .B(_01577_),
    .Y(_01647_)
  );
  XOR2X1 _08088_ (
    .A(_01574_),
    .B(_01577_),
    .Y(_01648_)
  );
  XNOR2X1 _08089_ (
    .A(_01646_),
    .B(_01647_),
    .Y(_01649_)
  );
  NAND2X1 _08090_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01646_),
    .Y(_01650_)
  );
  NAND2X1 _08091_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01638_),
    .Y(_01651_)
  );
  AOI21X1 _08092_ (
    .A(execution_unit_0.alu_0.alu_swpb_8_ ),
    .B(execution_unit_0.alu_0.inst_so_1_ ),
    .C(_01621_),
    .Y(_01652_)
  );
  OAI21X1 _08093_ (
    .A(_01375_),
    .B(_01645_),
    .C(_01652_),
    .Y(_01653_)
  );
  AOI22X1 _08094_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_8_ ),
    .C(_01415_),
    .D(_01637_),
    .Y(_01654_)
  );
  NAND3X1 _08095_ (
    .A(_01650_),
    .B(_01651_),
    .C(_01654_),
    .Y(_01655_)
  );
  OAI21X1 _08096_ (
    .A(_01653_),
    .B(_01655_),
    .C(_01386_),
    .Y(_01656_)
  );
  AOI22X1 _08097_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01649_),
    .C(_01656_),
    .D(_01504_),
    .Y(_01657_)
  );
  INVX1 _08098_ (
    .A(_01657_),
    .Y(_01658_)
  );
  NOR2X1 _08099_ (
    .A(_01613_),
    .B(_01644_),
    .Y(_01659_)
  );
  XNOR2X1 _08100_ (
    .A(_01613_),
    .B(_01644_),
    .Y(_01660_)
  );
  OAI21X1 _08101_ (
    .A(_01386_),
    .B(_01660_),
    .C(_01658_),
    .Y(execution_unit_0.alu_0.alu_out_8_ )
  );
  XNOR2X1 _08102_ (
    .A(execution_unit_0.alu_0.alu_shift_8_ ),
    .B(_01388_),
    .Y(_01661_)
  );
  NOR2X1 _08103_ (
    .A(_01634_),
    .B(_01661_),
    .Y(_01662_)
  );
  AND2X1 _08104_ (
    .A(execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01662_),
    .Y(_01663_)
  );
  NAND2X1 _08105_ (
    .A(execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01662_),
    .Y(_01664_)
  );
  NOR2X1 _08106_ (
    .A(_01401_),
    .B(_01664_),
    .Y(_01665_)
  );
  AOI21X1 _08107_ (
    .A(execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01635_),
    .C(_01662_),
    .Y(_01666_)
  );
  AOI22X1 _08108_ (
    .A(execution_unit_0.alu_0.op_dst_9_ ),
    .B(_01635_),
    .C(_01662_),
    .D(_01400_),
    .Y(_01667_)
  );
  NOR2X1 _08109_ (
    .A(_01665_),
    .B(_01667_),
    .Y(_01668_)
  );
  OAI21X1 _08110_ (
    .A(_01401_),
    .B(_01639_),
    .C(_01643_),
    .Y(_01669_)
  );
  XOR2X1 _08111_ (
    .A(_01668_),
    .B(_01669_),
    .Y(dbg_0.UNUSED_eu_mab_9_ )
  );
  NOR2X1 _08112_ (
    .A(_01659_),
    .B(dbg_0.UNUSED_eu_mab_9_ ),
    .Y(_01670_)
  );
  NAND2X1 _08113_ (
    .A(_01659_),
    .B(dbg_0.UNUSED_eu_mab_9_ ),
    .Y(_01671_)
  );
  OAI21X1 _08114_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01385_),
    .C(_01671_),
    .Y(_01672_)
  );
  NOR2X1 _08115_ (
    .A(_01663_),
    .B(_01666_),
    .Y(_01673_)
  );
  AOI21X1 _08116_ (
    .A(_01646_),
    .B(_01647_),
    .C(_01638_),
    .Y(_01674_)
  );
  OAI21X1 _08117_ (
    .A(_01645_),
    .B(_01648_),
    .C(_01639_),
    .Y(_01675_)
  );
  XNOR2X1 _08118_ (
    .A(_01673_),
    .B(_01674_),
    .Y(_01676_)
  );
  XNOR2X1 _08119_ (
    .A(execution_unit_0.alu_0.alu_shift_10_ ),
    .B(_01388_),
    .Y(_01677_)
  );
  NOR2X1 _08120_ (
    .A(_01634_),
    .B(_01677_),
    .Y(_01678_)
  );
  AND2X1 _08121_ (
    .A(execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01678_),
    .Y(_01679_)
  );
  NAND2X1 _08122_ (
    .A(execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01678_),
    .Y(_01680_)
  );
  AOI21X1 _08123_ (
    .A(execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01635_),
    .C(_01678_),
    .Y(_01681_)
  );
  NOR2X1 _08124_ (
    .A(_01679_),
    .B(_01681_),
    .Y(_01682_)
  );
  XNOR2X1 _08125_ (
    .A(execution_unit_0.alu_0.alu_shift_9_ ),
    .B(_01388_),
    .Y(_01683_)
  );
  NOR2X1 _08126_ (
    .A(_01634_),
    .B(_01683_),
    .Y(_01684_)
  );
  OAI21X1 _08127_ (
    .A(_01919_),
    .B(_01383_),
    .C(execution_unit_0.alu_0.op_dst_10_ ),
    .Y(_01685_)
  );
  NOR2X1 _08128_ (
    .A(_01683_),
    .B(_01685_),
    .Y(_01686_)
  );
  INVX1 _08129_ (
    .A(_01686_),
    .Y(_01687_)
  );
  AOI21X1 _08130_ (
    .A(_01673_),
    .B(_01675_),
    .C(_01663_),
    .Y(_01688_)
  );
  OAI21X1 _08131_ (
    .A(_01666_),
    .B(_01674_),
    .C(_01664_),
    .Y(_01689_)
  );
  AOI21X1 _08132_ (
    .A(execution_unit_0.alu_0.op_dst_10_ ),
    .B(_01635_),
    .C(_01684_),
    .Y(_01690_)
  );
  NOR2X1 _08133_ (
    .A(_01686_),
    .B(_01690_),
    .Y(_01691_)
  );
  AOI21X1 _08134_ (
    .A(_01689_),
    .B(_01691_),
    .C(_01686_),
    .Y(_01692_)
  );
  OAI21X1 _08135_ (
    .A(_01688_),
    .B(_01690_),
    .C(_01687_),
    .Y(_01693_)
  );
  AOI21X1 _08136_ (
    .A(_01682_),
    .B(_01693_),
    .C(_01679_),
    .Y(_01694_)
  );
  OAI21X1 _08137_ (
    .A(_01681_),
    .B(_01692_),
    .C(_01680_),
    .Y(_01695_)
  );
  XNOR2X1 _08138_ (
    .A(_01682_),
    .B(_01692_),
    .Y(_01696_)
  );
  XNOR2X1 _08139_ (
    .A(_01682_),
    .B(_01693_),
    .Y(_01697_)
  );
  XNOR2X1 _08140_ (
    .A(_01688_),
    .B(_01691_),
    .Y(_01698_)
  );
  NOR2X1 _08141_ (
    .A(_01676_),
    .B(_01698_),
    .Y(_01699_)
  );
  OR2X1 _08142_ (
    .A(_01676_),
    .B(_01698_),
    .Y(_01700_)
  );
  AOI21X1 _08143_ (
    .A(_01696_),
    .B(_01700_),
    .C(_01695_),
    .Y(_01701_)
  );
  OAI21X1 _08144_ (
    .A(_01697_),
    .B(_01699_),
    .C(_01694_),
    .Y(_01702_)
  );
  NOR2X1 _08145_ (
    .A(_01676_),
    .B(_01701_),
    .Y(_01703_)
  );
  XNOR2X1 _08146_ (
    .A(_01676_),
    .B(_01702_),
    .Y(_01704_)
  );
  NAND2X1 _08147_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01673_),
    .Y(_01705_)
  );
  NAND2X1 _08148_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01663_),
    .Y(_01706_)
  );
  AOI21X1 _08149_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_0_ ),
    .C(_01621_),
    .Y(_01707_)
  );
  OAI21X1 _08150_ (
    .A(_01375_),
    .B(_01666_),
    .C(_01707_),
    .Y(_01708_)
  );
  AOI22X1 _08151_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_9_ ),
    .C(_01415_),
    .D(_01662_),
    .Y(_01709_)
  );
  NAND3X1 _08152_ (
    .A(_01705_),
    .B(_01706_),
    .C(_01709_),
    .Y(_01710_)
  );
  OAI21X1 _08153_ (
    .A(_01708_),
    .B(_01710_),
    .C(_01386_),
    .Y(_01711_)
  );
  AOI22X1 _08154_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01704_),
    .C(_01711_),
    .D(_01504_),
    .Y(_01712_)
  );
  INVX1 _08155_ (
    .A(_01712_),
    .Y(_01713_)
  );
  OAI21X1 _08156_ (
    .A(_01670_),
    .B(_01672_),
    .C(_01713_),
    .Y(execution_unit_0.alu_0.alu_out_9_ )
  );
  NOR2X1 _08157_ (
    .A(_01640_),
    .B(_01666_),
    .Y(_01714_)
  );
  NOR2X1 _08158_ (
    .A(_01665_),
    .B(_01714_),
    .Y(_01715_)
  );
  OAI21X1 _08159_ (
    .A(_01643_),
    .B(_01667_),
    .C(_01715_),
    .Y(_01716_)
  );
  NAND2X1 _08160_ (
    .A(_01400_),
    .B(_01684_),
    .Y(_01717_)
  );
  NAND2X1 _08161_ (
    .A(_01400_),
    .B(_01686_),
    .Y(_01718_)
  );
  AOI22X1 _08162_ (
    .A(_01400_),
    .B(_01686_),
    .C(_01717_),
    .D(_01685_),
    .Y(_01719_)
  );
  NAND2X1 _08163_ (
    .A(_01716_),
    .B(_01719_),
    .Y(_01720_)
  );
  XNOR2X1 _08164_ (
    .A(_01716_),
    .B(_01719_),
    .Y(_01721_)
  );
  INVX1 _08165_ (
    .A(_01721_),
    .Y(dbg_0.UNUSED_eu_mab_10_ )
  );
  NAND2X1 _08166_ (
    .A(_01671_),
    .B(_01721_),
    .Y(_01722_)
  );
  OR2X1 _08167_ (
    .A(_01671_),
    .B(_01721_),
    .Y(_01723_)
  );
  NAND2X1 _08168_ (
    .A(_01722_),
    .B(_01723_),
    .Y(_01724_)
  );
  AOI21X1 _08169_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_1_ ),
    .C(_01621_),
    .Y(_01725_)
  );
  AOI22X1 _08170_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_10_ ),
    .C(_01415_),
    .D(_01684_),
    .Y(_01726_)
  );
  OAI21X1 _08171_ (
    .A(_01376_),
    .B(_01687_),
    .C(_01726_),
    .Y(_01727_)
  );
  OAI21X1 _08172_ (
    .A(_01375_),
    .B(_01690_),
    .C(_01725_),
    .Y(_01728_)
  );
  NOR2X1 _08173_ (
    .A(_01727_),
    .B(_01728_),
    .Y(_01729_)
  );
  AOI21X1 _08174_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01691_),
    .C(_01387_),
    .Y(_01730_)
  );
  NAND2X1 _08175_ (
    .A(_01729_),
    .B(_01730_),
    .Y(_01731_)
  );
  OAI21X1 _08176_ (
    .A(_01379_),
    .B(_01387_),
    .C(_01731_),
    .Y(_01732_)
  );
  AOI21X1 _08177_ (
    .A(_01698_),
    .B(_01703_),
    .C(_01379_),
    .Y(_01733_)
  );
  OAI21X1 _08178_ (
    .A(_01698_),
    .B(_01703_),
    .C(_01733_),
    .Y(_01734_)
  );
  AOI22X1 _08179_ (
    .A(_01387_),
    .B(_01724_),
    .C(_01732_),
    .D(_01734_),
    .Y(execution_unit_0.alu_0.alu_out_10_ )
  );
  OAI21X1 _08180_ (
    .A(_01401_),
    .B(_01687_),
    .C(_01720_),
    .Y(_01735_)
  );
  NOR2X1 _08181_ (
    .A(_01401_),
    .B(_01680_),
    .Y(_01736_)
  );
  AOI22X1 _08182_ (
    .A(execution_unit_0.alu_0.op_dst_11_ ),
    .B(_01635_),
    .C(_01678_),
    .D(_01400_),
    .Y(_01737_)
  );
  NOR2X1 _08183_ (
    .A(_01736_),
    .B(_01737_),
    .Y(_01738_)
  );
  XNOR2X1 _08184_ (
    .A(_01735_),
    .B(_01738_),
    .Y(_01739_)
  );
  INVX1 _08185_ (
    .A(_01739_),
    .Y(dbg_0.UNUSED_eu_mab_11_ )
  );
  NOR2X1 _08186_ (
    .A(_01723_),
    .B(_01739_),
    .Y(_01740_)
  );
  XNOR2X1 _08187_ (
    .A(_01723_),
    .B(_01739_),
    .Y(_01741_)
  );
  AOI21X1 _08188_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_2_ ),
    .C(_01621_),
    .Y(_01742_)
  );
  AOI22X1 _08189_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_11_ ),
    .C(_01415_),
    .D(_01678_),
    .Y(_01743_)
  );
  OAI21X1 _08190_ (
    .A(_01376_),
    .B(_01680_),
    .C(_01743_),
    .Y(_01744_)
  );
  OAI21X1 _08191_ (
    .A(_01375_),
    .B(_01681_),
    .C(_01742_),
    .Y(_01745_)
  );
  NOR2X1 _08192_ (
    .A(_01744_),
    .B(_01745_),
    .Y(_01746_)
  );
  AOI21X1 _08193_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01682_),
    .C(_01387_),
    .Y(_01747_)
  );
  NAND2X1 _08194_ (
    .A(_01746_),
    .B(_01747_),
    .Y(_01748_)
  );
  OAI21X1 _08195_ (
    .A(_01694_),
    .B(_01699_),
    .C(_01697_),
    .Y(_01749_)
  );
  AOI21X1 _08196_ (
    .A(_01696_),
    .B(_01700_),
    .C(_01379_),
    .Y(_01750_)
  );
  AOI22X1 _08197_ (
    .A(_01504_),
    .B(_01748_),
    .C(_01749_),
    .D(_01750_),
    .Y(_01751_)
  );
  AOI21X1 _08198_ (
    .A(_01387_),
    .B(_01741_),
    .C(_01751_),
    .Y(execution_unit_0.alu_0.alu_out_11_ )
  );
  AOI21X1 _08199_ (
    .A(_01718_),
    .B(_01720_),
    .C(_01737_),
    .Y(_01752_)
  );
  OR2X1 _08200_ (
    .A(_01736_),
    .B(_01752_),
    .Y(_01753_)
  );
  OAI21X1 _08201_ (
    .A(execution_unit_0.alu_0.alu_shift_11_ ),
    .B(_01388_),
    .C(_01635_),
    .Y(_01754_)
  );
  AOI21X1 _08202_ (
    .A(execution_unit_0.alu_0.alu_shift_11_ ),
    .B(_01388_),
    .C(_01754_),
    .Y(_01755_)
  );
  AND2X1 _08203_ (
    .A(execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01755_),
    .Y(_01756_)
  );
  NAND2X1 _08204_ (
    .A(execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01755_),
    .Y(_01757_)
  );
  AOI22X1 _08205_ (
    .A(execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01635_),
    .C(_01755_),
    .D(_01400_),
    .Y(_01758_)
  );
  AOI21X1 _08206_ (
    .A(_01400_),
    .B(_01756_),
    .C(_01758_),
    .Y(_01759_)
  );
  XOR2X1 _08207_ (
    .A(_01753_),
    .B(_01759_),
    .Y(dbg_0.UNUSED_eu_mab_12_ )
  );
  AND2X1 _08208_ (
    .A(_01740_),
    .B(dbg_0.UNUSED_eu_mab_12_ ),
    .Y(_01760_)
  );
  OAI21X1 _08209_ (
    .A(_01740_),
    .B(dbg_0.UNUSED_eu_mab_12_ ),
    .C(_01387_),
    .Y(_01761_)
  );
  OR2X1 _08210_ (
    .A(_01760_),
    .B(_01761_),
    .Y(_01762_)
  );
  AOI21X1 _08211_ (
    .A(execution_unit_0.alu_0.op_dst_12_ ),
    .B(_01635_),
    .C(_01755_),
    .Y(_01763_)
  );
  NOR2X1 _08212_ (
    .A(_01756_),
    .B(_01763_),
    .Y(_01764_)
  );
  INVX1 _08213_ (
    .A(_01764_),
    .Y(_01765_)
  );
  NOR3X1 _08214_ (
    .A(_01694_),
    .B(_01697_),
    .C(_01699_),
    .Y(_01766_)
  );
  NAND3X1 _08215_ (
    .A(_01695_),
    .B(_01696_),
    .C(_01700_),
    .Y(_01767_)
  );
  NOR3X1 _08216_ (
    .A(_01701_),
    .B(_01765_),
    .C(_01766_),
    .Y(_01768_)
  );
  NAND3X1 _08217_ (
    .A(_01702_),
    .B(_01764_),
    .C(_01767_),
    .Y(_01769_)
  );
  OAI21X1 _08218_ (
    .A(_01701_),
    .B(_01766_),
    .C(_01765_),
    .Y(_01770_)
  );
  AND2X1 _08219_ (
    .A(_01769_),
    .B(_01770_),
    .Y(_01771_)
  );
  NAND2X1 _08220_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01764_),
    .Y(_01772_)
  );
  NAND2X1 _08221_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01756_),
    .Y(_01773_)
  );
  AOI21X1 _08222_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_3_ ),
    .C(_01621_),
    .Y(_01774_)
  );
  OAI21X1 _08223_ (
    .A(_01375_),
    .B(_01763_),
    .C(_01774_),
    .Y(_01775_)
  );
  AOI22X1 _08224_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_12_ ),
    .C(_01415_),
    .D(_01755_),
    .Y(_01776_)
  );
  NAND3X1 _08225_ (
    .A(_01772_),
    .B(_01773_),
    .C(_01776_),
    .Y(_01777_)
  );
  OAI21X1 _08226_ (
    .A(_01775_),
    .B(_01777_),
    .C(_01386_),
    .Y(_01778_)
  );
  OAI21X1 _08227_ (
    .A(_01379_),
    .B(_01387_),
    .C(_01778_),
    .Y(_01779_)
  );
  OAI21X1 _08228_ (
    .A(_01379_),
    .B(_01771_),
    .C(_01779_),
    .Y(_01780_)
  );
  OAI21X1 _08229_ (
    .A(_01760_),
    .B(_01761_),
    .C(_01780_),
    .Y(execution_unit_0.alu_0.alu_out_12_ )
  );
  XNOR2X1 _08230_ (
    .A(execution_unit_0.alu_0.alu_shift_12_ ),
    .B(_01388_),
    .Y(_01781_)
  );
  NOR2X1 _08231_ (
    .A(_01634_),
    .B(_01781_),
    .Y(_01782_)
  );
  AND2X1 _08232_ (
    .A(execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01782_),
    .Y(_01783_)
  );
  NAND2X1 _08233_ (
    .A(execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01782_),
    .Y(_01784_)
  );
  AOI21X1 _08234_ (
    .A(execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01635_),
    .C(_01782_),
    .Y(_01785_)
  );
  AOI22X1 _08235_ (
    .A(execution_unit_0.alu_0.op_dst_13_ ),
    .B(_01635_),
    .C(_01782_),
    .D(_01400_),
    .Y(_01786_)
  );
  AOI21X1 _08236_ (
    .A(_01400_),
    .B(_01783_),
    .C(_01786_),
    .Y(_01787_)
  );
  AOI22X1 _08237_ (
    .A(_01400_),
    .B(_01756_),
    .C(_01759_),
    .D(_01753_),
    .Y(_01788_)
  );
  XNOR2X1 _08238_ (
    .A(_01787_),
    .B(_01788_),
    .Y(dbg_0.UNUSED_eu_mab_13_ )
  );
  NOR2X1 _08239_ (
    .A(_01760_),
    .B(dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_01789_)
  );
  NAND2X1 _08240_ (
    .A(_01760_),
    .B(dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_01790_)
  );
  OAI21X1 _08241_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .B(_01385_),
    .C(_01790_),
    .Y(_01791_)
  );
  NOR2X1 _08242_ (
    .A(_01789_),
    .B(_01791_),
    .Y(_01792_)
  );
  NOR2X1 _08243_ (
    .A(_01783_),
    .B(_01785_),
    .Y(_01793_)
  );
  INVX1 _08244_ (
    .A(_01793_),
    .Y(_01794_)
  );
  NAND2X1 _08245_ (
    .A(_01757_),
    .B(_01769_),
    .Y(_01795_)
  );
  AOI21X1 _08246_ (
    .A(_01757_),
    .B(_01769_),
    .C(_01794_),
    .Y(_01796_)
  );
  OAI21X1 _08247_ (
    .A(_01756_),
    .B(_01768_),
    .C(_01793_),
    .Y(_01797_)
  );
  XNOR2X1 _08248_ (
    .A(_01794_),
    .B(_01795_),
    .Y(_01798_)
  );
  XNOR2X1 _08249_ (
    .A(_01793_),
    .B(_01795_),
    .Y(_01799_)
  );
  XNOR2X1 _08250_ (
    .A(execution_unit_0.alu_0.alu_shift_14_ ),
    .B(_01388_),
    .Y(_01800_)
  );
  NOR2X1 _08251_ (
    .A(_01634_),
    .B(_01800_),
    .Y(_01801_)
  );
  INVX1 _08252_ (
    .A(_01801_),
    .Y(_01802_)
  );
  NOR2X1 _08253_ (
    .A(_01384_),
    .B(_01802_),
    .Y(_01803_)
  );
  NAND2X1 _08254_ (
    .A(execution_unit_0.alu_0.op_dst_15_ ),
    .B(_01801_),
    .Y(_01804_)
  );
  OAI21X1 _08255_ (
    .A(_01384_),
    .B(_01634_),
    .C(_01802_),
    .Y(_01805_)
  );
  XNOR2X1 _08256_ (
    .A(execution_unit_0.alu_0.alu_shift_13_ ),
    .B(_01388_),
    .Y(_01806_)
  );
  NOR2X1 _08257_ (
    .A(_01634_),
    .B(_01806_),
    .Y(_01807_)
  );
  OAI21X1 _08258_ (
    .A(_01919_),
    .B(_01383_),
    .C(execution_unit_0.alu_0.op_dst_14_ ),
    .Y(_01808_)
  );
  NOR2X1 _08259_ (
    .A(_01806_),
    .B(_01808_),
    .Y(_01809_)
  );
  NAND2X1 _08260_ (
    .A(execution_unit_0.alu_0.op_dst_14_ ),
    .B(_01807_),
    .Y(_01810_)
  );
  OAI21X1 _08261_ (
    .A(_01634_),
    .B(_01806_),
    .C(_01808_),
    .Y(_01811_)
  );
  AND2X1 _08262_ (
    .A(_01810_),
    .B(_01811_),
    .Y(_01812_)
  );
  OAI21X1 _08263_ (
    .A(_01806_),
    .B(_01808_),
    .C(_01811_),
    .Y(_01813_)
  );
  AOI21X1 _08264_ (
    .A(_01784_),
    .B(_01797_),
    .C(_01813_),
    .Y(_01814_)
  );
  OAI21X1 _08265_ (
    .A(_01783_),
    .B(_01796_),
    .C(_01812_),
    .Y(_01815_)
  );
  OAI21X1 _08266_ (
    .A(_01809_),
    .B(_01814_),
    .C(_01805_),
    .Y(_01816_)
  );
  AND2X1 _08267_ (
    .A(_01804_),
    .B(_01816_),
    .Y(_01817_)
  );
  OAI21X1 _08268_ (
    .A(_01384_),
    .B(_01802_),
    .C(_01816_),
    .Y(_01818_)
  );
  NOR3X1 _08269_ (
    .A(_01783_),
    .B(_01796_),
    .C(_01812_),
    .Y(_01819_)
  );
  NAND3X1 _08270_ (
    .A(_01784_),
    .B(_01797_),
    .C(_01813_),
    .Y(_01820_)
  );
  NAND2X1 _08271_ (
    .A(_01815_),
    .B(_01820_),
    .Y(_01821_)
  );
  AOI21X1 _08272_ (
    .A(_01815_),
    .B(_01820_),
    .C(_01798_),
    .Y(_01822_)
  );
  OAI21X1 _08273_ (
    .A(_01814_),
    .B(_01819_),
    .C(_01799_),
    .Y(_01823_)
  );
  AND2X1 _08274_ (
    .A(_01804_),
    .B(_01805_),
    .Y(_01824_)
  );
  OAI21X1 _08275_ (
    .A(_01384_),
    .B(_01802_),
    .C(_01805_),
    .Y(_01825_)
  );
  OAI21X1 _08276_ (
    .A(_01809_),
    .B(_01814_),
    .C(_01825_),
    .Y(_01826_)
  );
  NAND3X1 _08277_ (
    .A(_01810_),
    .B(_01815_),
    .C(_01824_),
    .Y(_01827_)
  );
  NAND3X1 _08278_ (
    .A(_01810_),
    .B(_01815_),
    .C(_01825_),
    .Y(_01828_)
  );
  OAI21X1 _08279_ (
    .A(_01809_),
    .B(_01814_),
    .C(_01824_),
    .Y(_01829_)
  );
  NAND2X1 _08280_ (
    .A(_01828_),
    .B(_01829_),
    .Y(_01830_)
  );
  AOI21X1 _08281_ (
    .A(_01826_),
    .B(_01827_),
    .C(_01822_),
    .Y(_01831_)
  );
  NAND3X1 _08282_ (
    .A(_01823_),
    .B(_01828_),
    .C(_01829_),
    .Y(_01832_)
  );
  AOI21X1 _08283_ (
    .A(_01817_),
    .B(_01832_),
    .C(_01798_),
    .Y(_01833_)
  );
  OAI21X1 _08284_ (
    .A(_01818_),
    .B(_01831_),
    .C(_01799_),
    .Y(_01834_)
  );
  NAND3X1 _08285_ (
    .A(_01798_),
    .B(_01817_),
    .C(_01830_),
    .Y(_01835_)
  );
  NAND3X1 _08286_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01834_),
    .C(_01835_),
    .Y(_01836_)
  );
  NAND2X1 _08287_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01793_),
    .Y(_01837_)
  );
  NAND2X1 _08288_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01783_),
    .Y(_01838_)
  );
  AOI21X1 _08289_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_4_ ),
    .C(_01621_),
    .Y(_01839_)
  );
  OAI21X1 _08290_ (
    .A(_01375_),
    .B(_01785_),
    .C(_01839_),
    .Y(_01840_)
  );
  AOI22X1 _08291_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_13_ ),
    .C(_01415_),
    .D(_01782_),
    .Y(_01841_)
  );
  NAND3X1 _08292_ (
    .A(_01837_),
    .B(_01838_),
    .C(_01841_),
    .Y(_01842_)
  );
  OAI21X1 _08293_ (
    .A(_01840_),
    .B(_01842_),
    .C(_01386_),
    .Y(_01843_)
  );
  OAI21X1 _08294_ (
    .A(_01379_),
    .B(_01387_),
    .C(_01843_),
    .Y(_01844_)
  );
  AOI21X1 _08295_ (
    .A(_01836_),
    .B(_01844_),
    .C(_01792_),
    .Y(_01845_)
  );
  INVX1 _08296_ (
    .A(_01845_),
    .Y(execution_unit_0.alu_0.alu_out_13_ )
  );
  NAND2X1 _08297_ (
    .A(_01400_),
    .B(_01807_),
    .Y(_01846_)
  );
  AOI22X1 _08298_ (
    .A(_01400_),
    .B(_01809_),
    .C(_01846_),
    .D(_01808_),
    .Y(_01847_)
  );
  OAI22X1 _08299_ (
    .A(_01401_),
    .B(_01784_),
    .C(_01786_),
    .D(_01788_),
    .Y(_01848_)
  );
  NAND2X1 _08300_ (
    .A(_01847_),
    .B(_01848_),
    .Y(_01849_)
  );
  XNOR2X1 _08301_ (
    .A(_01847_),
    .B(_01848_),
    .Y(_01850_)
  );
  INVX1 _08302_ (
    .A(_01850_),
    .Y(dbg_0.UNUSED_eu_mab_14_ )
  );
  AOI21X1 _08303_ (
    .A(_01818_),
    .B(_01822_),
    .C(_01379_),
    .Y(_01851_)
  );
  OAI21X1 _08304_ (
    .A(_01821_),
    .B(_01833_),
    .C(_01851_),
    .Y(_01852_)
  );
  NAND2X1 _08305_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01811_),
    .Y(_01853_)
  );
  AOI21X1 _08306_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_5_ ),
    .C(_01621_),
    .Y(_01854_)
  );
  AOI22X1 _08307_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.alu_shift_14_ ),
    .C(_01415_),
    .D(_01807_),
    .Y(_01855_)
  );
  OAI21X1 _08308_ (
    .A(_01376_),
    .B(_01810_),
    .C(_01855_),
    .Y(_01856_)
  );
  AOI21X1 _08309_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_01812_),
    .C(_01856_),
    .Y(_01857_)
  );
  NAND3X1 _08310_ (
    .A(_01853_),
    .B(_01854_),
    .C(_01857_),
    .Y(_01858_)
  );
  OAI21X1 _08311_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .B(_01858_),
    .C(_01386_),
    .Y(_01859_)
  );
  INVX1 _08312_ (
    .A(_01859_),
    .Y(_01860_)
  );
  OR2X1 _08313_ (
    .A(_01790_),
    .B(_01850_),
    .Y(_01861_)
  );
  AOI21X1 _08314_ (
    .A(_01790_),
    .B(_01850_),
    .C(_01386_),
    .Y(_01862_)
  );
  AND2X1 _08315_ (
    .A(_01861_),
    .B(_01862_),
    .Y(_01863_)
  );
  AOI21X1 _08316_ (
    .A(_01852_),
    .B(_01860_),
    .C(_01863_),
    .Y(_01864_)
  );
  INVX1 _08317_ (
    .A(_01864_),
    .Y(execution_unit_0.alu_0.alu_out_14_ )
  );
  OAI21X1 _08318_ (
    .A(_01401_),
    .B(_01810_),
    .C(_01849_),
    .Y(_01865_)
  );
  AOI22X1 _08319_ (
    .A(execution_unit_0.alu_0.op_dst_15_ ),
    .B(_01635_),
    .C(_01801_),
    .D(_01400_),
    .Y(_01866_)
  );
  AOI21X1 _08320_ (
    .A(_01400_),
    .B(_01803_),
    .C(_01866_),
    .Y(_01867_)
  );
  NAND2X1 _08321_ (
    .A(_01865_),
    .B(_01867_),
    .Y(_01868_)
  );
  XNOR2X1 _08322_ (
    .A(_01865_),
    .B(_01867_),
    .Y(_01869_)
  );
  INVX1 _08323_ (
    .A(_01869_),
    .Y(dbg_0.UNUSED_eu_mab_15_ )
  );
  NOR2X1 _08324_ (
    .A(_01861_),
    .B(_01869_),
    .Y(_01870_)
  );
  AND2X1 _08325_ (
    .A(_01861_),
    .B(_01869_),
    .Y(_01871_)
  );
  OAI21X1 _08326_ (
    .A(_01870_),
    .B(_01871_),
    .C(_01387_),
    .Y(_01872_)
  );
  NAND2X1 _08327_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(execution_unit_0.alu_0.alu_shift_6_ ),
    .Y(_01873_)
  );
  AOI22X1 _08328_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(_01617_),
    .C(_01801_),
    .D(_01415_),
    .Y(_01874_)
  );
  AOI21X1 _08329_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_01803_),
    .C(_01621_),
    .Y(_01875_)
  );
  NAND2X1 _08330_ (
    .A(_01873_),
    .B(_01874_),
    .Y(_01876_)
  );
  AOI21X1 _08331_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_01805_),
    .C(_01876_),
    .Y(_01877_)
  );
  NAND2X1 _08332_ (
    .A(_01875_),
    .B(_01877_),
    .Y(_01878_)
  );
  OAI21X1 _08333_ (
    .A(_01374_),
    .B(_01825_),
    .C(_01386_),
    .Y(_01879_)
  );
  OAI21X1 _08334_ (
    .A(_01878_),
    .B(_01879_),
    .C(_01504_),
    .Y(_01880_)
  );
  AOI22X1 _08335_ (
    .A(_01818_),
    .B(_01823_),
    .C(_01828_),
    .D(_01829_),
    .Y(_01881_)
  );
  OAI21X1 _08336_ (
    .A(_01822_),
    .B(_01830_),
    .C(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_01882_)
  );
  OAI21X1 _08337_ (
    .A(_01881_),
    .B(_01882_),
    .C(_01880_),
    .Y(_01883_)
  );
  NAND2X1 _08338_ (
    .A(_01872_),
    .B(_01883_),
    .Y(_01884_)
  );
  INVX1 _08339_ (
    .A(_01884_),
    .Y(execution_unit_0.alu_0.alu_out_15_ )
  );
  NAND2X1 _08340_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_01885_)
  );
  OAI21X1 _08341_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01884_),
    .C(_01885_),
    .Y(execution_unit_0.alu_0.N )
  );
  OR2X1 _08342_ (
    .A(execution_unit_0.alu_0.alu_out_8_ ),
    .B(execution_unit_0.alu_0.alu_out_11_ ),
    .Y(_01886_)
  );
  NOR3X1 _08343_ (
    .A(execution_unit_0.alu_0.alu_out_9_ ),
    .B(execution_unit_0.alu_0.alu_out_10_ ),
    .C(_01886_),
    .Y(_01887_)
  );
  NAND3X1 _08344_ (
    .A(_01762_),
    .B(_01780_),
    .C(_01887_),
    .Y(_01888_)
  );
  AOI21X1 _08345_ (
    .A(_01872_),
    .B(_01883_),
    .C(_01888_),
    .Y(_01889_)
  );
  NAND3X1 _08346_ (
    .A(_01845_),
    .B(_01864_),
    .C(_01889_),
    .Y(_01890_)
  );
  NOR2X1 _08347_ (
    .A(execution_unit_0.alu_0.alu_out_0_ ),
    .B(execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_01891_)
  );
  NAND2X1 _08348_ (
    .A(_01478_),
    .B(_01891_),
    .Y(_01892_)
  );
  NOR2X1 _08349_ (
    .A(execution_unit_0.alu_0.alu_out_2_ ),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_01893_)
  );
  NOR2X1 _08350_ (
    .A(execution_unit_0.alu_0.alu_out_4_ ),
    .B(_01892_),
    .Y(_01894_)
  );
  NAND2X1 _08351_ (
    .A(_01893_),
    .B(_01894_),
    .Y(_01895_)
  );
  OR2X1 _08352_ (
    .A(execution_unit_0.alu_0.alu_out_5_ ),
    .B(_01895_),
    .Y(_01896_)
  );
  OR2X1 _08353_ (
    .A(execution_unit_0.alu_0.alu_out_6_ ),
    .B(_01896_),
    .Y(_01897_)
  );
  AOI21X1 _08354_ (
    .A(_01383_),
    .B(_01890_),
    .C(_01897_),
    .Y(execution_unit_0.alu_0.Z )
  );
  NAND2X1 _08355_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(_01390_),
    .Y(_01898_)
  );
  OR2X1 _08356_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_01899_)
  );
  AND2X1 _08357_ (
    .A(execution_unit_0.alu_0.Z ),
    .B(_01899_),
    .Y(_01900_)
  );
  OAI21X1 _08358_ (
    .A(_01401_),
    .B(_01804_),
    .C(_01868_),
    .Y(_01901_)
  );
  OAI21X1 _08359_ (
    .A(_01870_),
    .B(_01901_),
    .C(_01387_),
    .Y(_01902_)
  );
  AOI21X1 _08360_ (
    .A(_01817_),
    .B(_01832_),
    .C(_01504_),
    .Y(_01903_)
  );
  OAI21X1 _08361_ (
    .A(_01817_),
    .B(_01832_),
    .C(_01903_),
    .Y(_01904_)
  );
  AOI21X1 _08362_ (
    .A(_01902_),
    .B(_01904_),
    .C(execution_unit_0.alu_0.inst_bw ),
    .Y(_01905_)
  );
  AND2X1 _08363_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(execution_unit_0.alu_0.alu_out_8_ ),
    .Y(_01906_)
  );
  OR2X1 _08364_ (
    .A(_01905_),
    .B(_01906_),
    .Y(_01907_)
  );
  OAI21X1 _08365_ (
    .A(_01899_),
    .B(_01907_),
    .C(_01377_),
    .Y(_01908_)
  );
  OAI21X1 _08366_ (
    .A(_01900_),
    .B(_01908_),
    .C(_01898_),
    .Y(execution_unit_0.alu_0.alu_stat_0_ )
  );
  OAI21X1 _08367_ (
    .A(execution_unit_0.alu_0.op_dst_7_ ),
    .B(_01566_),
    .C(execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_01909_)
  );
  OAI21X1 _08368_ (
    .A(_01567_),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .C(_01909_),
    .Y(_01910_)
  );
  NAND2X1 _08369_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01910_),
    .Y(_01911_)
  );
  NAND2X1 _08370_ (
    .A(_01803_),
    .B(_01884_),
    .Y(_01912_)
  );
  OAI21X1 _08371_ (
    .A(_01805_),
    .B(_01884_),
    .C(_01912_),
    .Y(_01913_)
  );
  OAI21X1 _08372_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01913_),
    .C(_01911_),
    .Y(_01914_)
  );
  AOI21X1 _08373_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01567_),
    .C(_01374_),
    .Y(_01915_)
  );
  OAI21X1 _08374_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_01804_),
    .C(_01915_),
    .Y(_01916_)
  );
  NOR2X1 _08375_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_01917_)
  );
  NAND2X1 _08376_ (
    .A(_01916_),
    .B(_01917_),
    .Y(_01918_)
  );
  AOI21X1 _08377_ (
    .A(_01374_),
    .B(_01914_),
    .C(_01918_),
    .Y(execution_unit_0.alu_0.alu_stat_3_ )
  );
  AND2X1 _08378_ (
    .A(execution_unit_0.alu_0.exec_cycle ),
    .B(execution_unit_0.alu_0.inst_alu_9_ ),
    .Y(execution_unit_0.alu_0.alu_stat_wr_0_ )
  );
  INVX1 _08379_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .Y(_02949_)
  );
  INVX1 _08380_ (
    .A(execution_unit_0.reg_sr_clr ),
    .Y(_02950_)
  );
  INVX1 _08381_ (
    .A(execution_unit_0.inst_src_1_ ),
    .Y(_02951_)
  );
  INVX1 _08382_ (
    .A(execution_unit_0.register_file_0.r9_0_ ),
    .Y(_02952_)
  );
  INVX1 _08383_ (
    .A(execution_unit_0.register_file_0.r10_0_ ),
    .Y(_02953_)
  );
  INVX1 _08384_ (
    .A(execution_unit_0.register_file_0.r15_0_ ),
    .Y(_02954_)
  );
  INVX1 _08385_ (
    .A(execution_unit_0.alu_0.alu_out_0_ ),
    .Y(_02955_)
  );
  INVX1 _08386_ (
    .A(execution_unit_0.alu_0.alu_out_1_ ),
    .Y(_02956_)
  );
  INVX1 _08387_ (
    .A(execution_unit_0.register_file_0.r1_2_ ),
    .Y(_02957_)
  );
  INVX1 _08388_ (
    .A(execution_unit_0.register_file_0.r15_2_ ),
    .Y(_02958_)
  );
  INVX1 _08389_ (
    .A(execution_unit_0.alu_0.alu_out_2_ ),
    .Y(_02959_)
  );
  INVX1 _08390_ (
    .A(execution_unit_0.register_file_0.r10_3_ ),
    .Y(_02960_)
  );
  INVX1 _08391_ (
    .A(execution_unit_0.register_file_0.r1_3_ ),
    .Y(_02961_)
  );
  INVX1 _08392_ (
    .A(execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_02962_)
  );
  INVX1 _08393_ (
    .A(execution_unit_0.register_file_0.r2_4_ ),
    .Y(_02963_)
  );
  INVX1 _08394_ (
    .A(execution_unit_0.register_file_0.r1_4_ ),
    .Y(_02964_)
  );
  INVX1 _08395_ (
    .A(execution_unit_0.alu_0.alu_out_4_ ),
    .Y(_02965_)
  );
  INVX1 _08396_ (
    .A(execution_unit_0.alu_0.alu_out_5_ ),
    .Y(_02966_)
  );
  INVX1 _08397_ (
    .A(execution_unit_0.alu_0.alu_out_6_ ),
    .Y(_02967_)
  );
  INVX1 _08398_ (
    .A(execution_unit_0.alu_0.alu_out_7_ ),
    .Y(_02968_)
  );
  INVX1 _08399_ (
    .A(execution_unit_0.register_file_0.r1_8_ ),
    .Y(_02969_)
  );
  INVX1 _08400_ (
    .A(execution_unit_0.register_file_0.r1_11_ ),
    .Y(_02970_)
  );
  INVX1 _08401_ (
    .A(execution_unit_0.register_file_0.r1_13_ ),
    .Y(_02971_)
  );
  INVX1 _08402_ (
    .A(execution_unit_0.register_file_0.r9_14_ ),
    .Y(_02972_)
  );
  INVX1 _08403_ (
    .A(execution_unit_0.register_file_0.r1_14_ ),
    .Y(_02973_)
  );
  INVX1 _08404_ (
    .A(execution_unit_0.register_file_0.r15_15_ ),
    .Y(_02974_)
  );
  INVX1 _08405_ (
    .A(execution_unit_0.register_file_0.r1_15_ ),
    .Y(_02975_)
  );
  INVX1 _08406_ (
    .A(execution_unit_0.inst_dest_9_ ),
    .Y(_02976_)
  );
  INVX1 _08407_ (
    .A(execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_02977_)
  );
  INVX1 _08408_ (
    .A(execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_02978_)
  );
  INVX1 _08409_ (
    .A(execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_02979_)
  );
  INVX1 _08410_ (
    .A(execution_unit_0.alu_0.alu_stat_wr_0_ ),
    .Y(_02980_)
  );
  INVX1 _08411_ (
    .A(execution_unit_0.reg_sp_wr ),
    .Y(_02981_)
  );
  INVX1 _08412_ (
    .A(_00162_),
    .Y(_02152_)
  );
  NAND2X1 _08413_ (
    .A(execution_unit_0.alu_0.alu_out_8_ ),
    .B(_02949_),
    .Y(_02982_)
  );
  INVX1 _08414_ (
    .A(_02982_),
    .Y(execution_unit_0.pc_sw_8_ )
  );
  NAND2X1 _08415_ (
    .A(_02949_),
    .B(execution_unit_0.alu_0.alu_out_9_ ),
    .Y(_02983_)
  );
  INVX1 _08416_ (
    .A(_02983_),
    .Y(execution_unit_0.pc_sw_9_ )
  );
  NAND2X1 _08417_ (
    .A(_02949_),
    .B(execution_unit_0.alu_0.alu_out_10_ ),
    .Y(_02984_)
  );
  INVX1 _08418_ (
    .A(_02984_),
    .Y(execution_unit_0.pc_sw_10_ )
  );
  NAND2X1 _08419_ (
    .A(_02949_),
    .B(execution_unit_0.alu_0.alu_out_11_ ),
    .Y(_02985_)
  );
  INVX1 _08420_ (
    .A(_02985_),
    .Y(execution_unit_0.pc_sw_11_ )
  );
  NAND2X1 _08421_ (
    .A(_02949_),
    .B(execution_unit_0.alu_0.alu_out_12_ ),
    .Y(_02986_)
  );
  INVX1 _08422_ (
    .A(_02986_),
    .Y(execution_unit_0.pc_sw_12_ )
  );
  NAND2X1 _08423_ (
    .A(_02949_),
    .B(execution_unit_0.alu_0.alu_out_13_ ),
    .Y(_02987_)
  );
  INVX1 _08424_ (
    .A(_02987_),
    .Y(execution_unit_0.pc_sw_13_ )
  );
  NAND2X1 _08425_ (
    .A(_02949_),
    .B(execution_unit_0.alu_0.alu_out_14_ ),
    .Y(_02988_)
  );
  INVX1 _08426_ (
    .A(_02988_),
    .Y(execution_unit_0.pc_sw_14_ )
  );
  NAND2X1 _08427_ (
    .A(_02949_),
    .B(execution_unit_0.alu_0.alu_out_15_ ),
    .Y(_02989_)
  );
  INVX1 _08428_ (
    .A(_02989_),
    .Y(execution_unit_0.pc_sw_15_ )
  );
  AND2X1 _08429_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_13_ ),
    .Y(_02990_)
  );
  NAND3X1 _08430_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_13_ ),
    .C(execution_unit_0.register_file_0.r13_0_ ),
    .Y(_02991_)
  );
  AND2X1 _08431_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_10_ ),
    .Y(_02992_)
  );
  NAND2X1 _08432_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_10_ ),
    .Y(_02993_)
  );
  OAI21X1 _08433_ (
    .A(_02953_),
    .B(_02993_),
    .C(_02991_),
    .Y(_02994_)
  );
  AND2X1 _08434_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_7_ ),
    .Y(_02995_)
  );
  NAND3X1 _08435_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_7_ ),
    .C(execution_unit_0.register_file_0.r7_0_ ),
    .Y(_02996_)
  );
  AND2X1 _08436_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_14_ ),
    .Y(_02997_)
  );
  NAND3X1 _08437_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_14_ ),
    .C(execution_unit_0.register_file_0.r14_0_ ),
    .Y(_02998_)
  );
  OR2X1 _08438_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(execution_unit_0.inst_src_2_ ),
    .Y(_02999_)
  );
  OAI21X1 _08439_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(execution_unit_0.inst_src_2_ ),
    .C(execution_unit_0.alu_0.status_0_ ),
    .Y(_03000_)
  );
  NOR2X1 _08440_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02951_),
    .Y(_03001_)
  );
  NAND2X1 _08441_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_1_ ),
    .Y(_03002_)
  );
  NAND3X1 _08442_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_1_ ),
    .C(execution_unit_0.register_file_0.r1_0_ ),
    .Y(_03003_)
  );
  AND2X1 _08443_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_5_ ),
    .Y(_03004_)
  );
  AND2X1 _08444_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_3_ ),
    .Y(_03005_)
  );
  NAND3X1 _08445_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_3_ ),
    .C(execution_unit_0.register_file_0.r3_0_ ),
    .Y(_03006_)
  );
  AND2X1 _08446_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_4_ ),
    .Y(_03007_)
  );
  NAND3X1 _08447_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_4_ ),
    .C(execution_unit_0.register_file_0.r4_0_ ),
    .Y(_03008_)
  );
  AND2X1 _08448_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_11_ ),
    .Y(_03009_)
  );
  NAND3X1 _08449_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_11_ ),
    .C(execution_unit_0.register_file_0.r11_0_ ),
    .Y(_03010_)
  );
  AND2X1 _08450_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_12_ ),
    .Y(_03011_)
  );
  NAND3X1 _08451_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_12_ ),
    .C(execution_unit_0.register_file_0.r12_0_ ),
    .Y(_03012_)
  );
  AND2X1 _08452_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_6_ ),
    .Y(_03013_)
  );
  NAND3X1 _08453_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_6_ ),
    .C(execution_unit_0.register_file_0.r6_0_ ),
    .Y(_03014_)
  );
  AND2X1 _08454_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_0_ ),
    .Y(_03015_)
  );
  NAND3X1 _08455_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_0_ ),
    .C(dbg_0.UNUSED_pc_0_ ),
    .Y(_03016_)
  );
  AND2X1 _08456_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_9_ ),
    .Y(_03017_)
  );
  NAND2X1 _08457_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_9_ ),
    .Y(_03018_)
  );
  OAI21X1 _08458_ (
    .A(_02952_),
    .B(_03018_),
    .C(_03016_),
    .Y(_03019_)
  );
  AND2X1 _08459_ (
    .A(execution_unit_0.inst_src_15_ ),
    .B(_02950_),
    .Y(_03020_)
  );
  NAND2X1 _08460_ (
    .A(execution_unit_0.inst_src_15_ ),
    .B(_02950_),
    .Y(_03021_)
  );
  AND2X1 _08461_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_8_ ),
    .Y(_03022_)
  );
  NAND3X1 _08462_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_8_ ),
    .C(execution_unit_0.register_file_0.r8_0_ ),
    .Y(_03023_)
  );
  OAI21X1 _08463_ (
    .A(_02954_),
    .B(_03021_),
    .C(_03023_),
    .Y(_03024_)
  );
  NAND3X1 _08464_ (
    .A(_03000_),
    .B(_03003_),
    .C(_03008_),
    .Y(_03025_)
  );
  NAND3X1 _08465_ (
    .A(_02996_),
    .B(_02998_),
    .C(_03010_),
    .Y(_03026_)
  );
  NOR2X1 _08466_ (
    .A(_03025_),
    .B(_03026_),
    .Y(_03027_)
  );
  NOR3X1 _08467_ (
    .A(_02994_),
    .B(_03019_),
    .C(_03024_),
    .Y(_03028_)
  );
  NAND3X1 _08468_ (
    .A(_03006_),
    .B(_03012_),
    .C(_03014_),
    .Y(_03029_)
  );
  AOI21X1 _08469_ (
    .A(execution_unit_0.register_file_0.r5_0_ ),
    .B(_03004_),
    .C(_03029_),
    .Y(_03030_)
  );
  NAND3X1 _08470_ (
    .A(_03027_),
    .B(_03028_),
    .C(_03030_),
    .Y(execution_unit_0.reg_src_0_ )
  );
  AND2X1 _08471_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.reg_dest_wr ),
    .Y(_03031_)
  );
  NAND2X1 _08472_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.reg_dest_wr ),
    .Y(_03032_)
  );
  AND2X1 _08473_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03020_),
    .Y(_03033_)
  );
  NAND2X1 _08474_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03020_),
    .Y(_03034_)
  );
  OAI21X1 _08475_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02951_),
    .C(execution_unit_0.alu_0.inst_bw ),
    .Y(_03035_)
  );
  NOR2X1 _08476_ (
    .A(execution_unit_0.reg_src_0_ ),
    .B(_03035_),
    .Y(_03036_)
  );
  XOR2X1 _08477_ (
    .A(execution_unit_0.reg_src_0_ ),
    .B(_03035_),
    .Y(_03037_)
  );
  AOI21X1 _08478_ (
    .A(_03033_),
    .B(_03037_),
    .C(_03031_),
    .Y(_03038_)
  );
  OAI21X1 _08479_ (
    .A(execution_unit_0.register_file_0.r15_0_ ),
    .B(_03033_),
    .C(_03038_),
    .Y(_03039_)
  );
  OAI21X1 _08480_ (
    .A(_02955_),
    .B(_03032_),
    .C(_03039_),
    .Y(_02000_)
  );
  NAND3X1 _08481_ (
    .A(execution_unit_0.inst_src_15_ ),
    .B(_02950_),
    .C(execution_unit_0.register_file_0.r15_1_ ),
    .Y(_03040_)
  );
  OAI21X1 _08482_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(execution_unit_0.inst_src_2_ ),
    .C(execution_unit_0.alu_0.status_1_ ),
    .Y(_03041_)
  );
  NAND3X1 _08483_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_1_ ),
    .C(execution_unit_0.register_file_0.r1_1_ ),
    .Y(_03042_)
  );
  NAND3X1 _08484_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_8_ ),
    .C(execution_unit_0.register_file_0.r8_1_ ),
    .Y(_03043_)
  );
  NAND3X1 _08485_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_0_ ),
    .C(dbg_0.UNUSED_pc_1_ ),
    .Y(_03044_)
  );
  NAND3X1 _08486_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_10_ ),
    .C(execution_unit_0.register_file_0.r10_1_ ),
    .Y(_03045_)
  );
  NAND3X1 _08487_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_9_ ),
    .C(execution_unit_0.register_file_0.r9_1_ ),
    .Y(_03046_)
  );
  NAND3X1 _08488_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_14_ ),
    .C(execution_unit_0.register_file_0.r14_1_ ),
    .Y(_03047_)
  );
  NAND3X1 _08489_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_12_ ),
    .C(execution_unit_0.register_file_0.r12_1_ ),
    .Y(_03048_)
  );
  NAND3X1 _08490_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_6_ ),
    .C(execution_unit_0.register_file_0.r6_1_ ),
    .Y(_03049_)
  );
  NAND3X1 _08491_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_13_ ),
    .C(execution_unit_0.register_file_0.r13_1_ ),
    .Y(_03050_)
  );
  NAND3X1 _08492_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_4_ ),
    .C(execution_unit_0.register_file_0.r4_1_ ),
    .Y(_03051_)
  );
  AOI22X1 _08493_ (
    .A(execution_unit_0.register_file_0.r5_1_ ),
    .B(_03004_),
    .C(_03009_),
    .D(execution_unit_0.register_file_0.r11_1_ ),
    .Y(_03052_)
  );
  AOI22X1 _08494_ (
    .A(execution_unit_0.register_file_0.r7_1_ ),
    .B(_02995_),
    .C(_03005_),
    .D(execution_unit_0.register_file_0.r3_1_ ),
    .Y(_03053_)
  );
  AND2X1 _08495_ (
    .A(_03052_),
    .B(_03053_),
    .Y(_03054_)
  );
  NAND3X1 _08496_ (
    .A(_03040_),
    .B(_03046_),
    .C(_03050_),
    .Y(_03055_)
  );
  NAND3X1 _08497_ (
    .A(_03041_),
    .B(_03047_),
    .C(_03051_),
    .Y(_03056_)
  );
  NOR2X1 _08498_ (
    .A(_03055_),
    .B(_03056_),
    .Y(_03057_)
  );
  NAND3X1 _08499_ (
    .A(_03042_),
    .B(_03044_),
    .C(_03045_),
    .Y(_03058_)
  );
  NAND3X1 _08500_ (
    .A(_03043_),
    .B(_03048_),
    .C(_03049_),
    .Y(_03059_)
  );
  NOR2X1 _08501_ (
    .A(_03058_),
    .B(_03059_),
    .Y(_03060_)
  );
  NAND3X1 _08502_ (
    .A(_03054_),
    .B(_03057_),
    .C(_03060_),
    .Y(execution_unit_0.reg_src_1_ )
  );
  OAI21X1 _08503_ (
    .A(execution_unit_0.reg_src_0_ ),
    .B(_03035_),
    .C(execution_unit_0.reg_src_1_ ),
    .Y(_03061_)
  );
  XNOR2X1 _08504_ (
    .A(_03036_),
    .B(execution_unit_0.reg_src_1_ ),
    .Y(_03062_)
  );
  NOR2X1 _08505_ (
    .A(execution_unit_0.register_file_0.r15_1_ ),
    .B(_03033_),
    .Y(_03063_)
  );
  OAI21X1 _08506_ (
    .A(_03034_),
    .B(_03062_),
    .C(_03032_),
    .Y(_03064_)
  );
  OAI22X1 _08507_ (
    .A(_02956_),
    .B(_03032_),
    .C(_03063_),
    .D(_03064_),
    .Y(_02007_)
  );
  NAND3X1 _08508_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_5_ ),
    .C(execution_unit_0.register_file_0.r5_2_ ),
    .Y(_03065_)
  );
  NAND3X1 _08509_ (
    .A(_02950_),
    .B(execution_unit_0.inst_src_11_ ),
    .C(execution_unit_0.register_file_0.r11_2_ ),
    .Y(_03066_)
  );
  OAI21X1 _08510_ (
    .A(_02958_),
    .B(_03021_),
    .C(_03066_),
    .Y(_03067_)
  );
  AOI22X1 _08511_ (
    .A(execution_unit_0.register_file_0.r4_2_ ),
    .B(_03007_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_2_ ),
    .Y(_03068_)
  );
  AND2X1 _08512_ (
    .A(execution_unit_0.register_file_0.r14_2_ ),
    .B(_02997_),
    .Y(_03069_)
  );
  NAND2X1 _08513_ (
    .A(execution_unit_0.register_file_0.r12_2_ ),
    .B(_03011_),
    .Y(_03070_)
  );
  AOI22X1 _08514_ (
    .A(execution_unit_0.register_file_0.r3_2_ ),
    .B(_03005_),
    .C(_03015_),
    .D(dbg_0.UNUSED_pc_2_ ),
    .Y(_03071_)
  );
  OAI21X1 _08515_ (
    .A(_02957_),
    .B(_03002_),
    .C(_03065_),
    .Y(_03072_)
  );
  NOR3X1 _08516_ (
    .A(_03067_),
    .B(_03069_),
    .C(_03072_),
    .Y(_03073_)
  );
  NAND2X1 _08517_ (
    .A(_03070_),
    .B(_03071_),
    .Y(_03074_)
  );
  AOI22X1 _08518_ (
    .A(execution_unit_0.register_file_0.r10_2_ ),
    .B(_02992_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_2_ ),
    .Y(_03075_)
  );
  AOI22X1 _08519_ (
    .A(execution_unit_0.alu_0.status_2_ ),
    .B(_02999_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_2_ ),
    .Y(_03076_)
  );
  AND2X1 _08520_ (
    .A(_03075_),
    .B(_03076_),
    .Y(_03077_)
  );
  AOI22X1 _08521_ (
    .A(execution_unit_0.register_file_0.r13_2_ ),
    .B(_02990_),
    .C(_02995_),
    .D(execution_unit_0.register_file_0.r7_2_ ),
    .Y(_03078_)
  );
  AND2X1 _08522_ (
    .A(_03068_),
    .B(_03078_),
    .Y(_03079_)
  );
  NAND3X1 _08523_ (
    .A(_03073_),
    .B(_03077_),
    .C(_03079_),
    .Y(_03080_)
  );
  NOR2X1 _08524_ (
    .A(_03074_),
    .B(_03080_),
    .Y(_03081_)
  );
  INVX1 _08525_ (
    .A(_03081_),
    .Y(execution_unit_0.reg_src_2_ )
  );
  NOR2X1 _08526_ (
    .A(_03061_),
    .B(_03081_),
    .Y(_03082_)
  );
  XNOR2X1 _08527_ (
    .A(_03061_),
    .B(_03081_),
    .Y(_03083_)
  );
  AOI21X1 _08528_ (
    .A(_03033_),
    .B(_03083_),
    .C(_03031_),
    .Y(_03084_)
  );
  OAI21X1 _08529_ (
    .A(execution_unit_0.register_file_0.r15_2_ ),
    .B(_03033_),
    .C(_03084_),
    .Y(_03085_)
  );
  OAI21X1 _08530_ (
    .A(_02959_),
    .B(_03032_),
    .C(_03085_),
    .Y(_02008_)
  );
  OAI21X1 _08531_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(execution_unit_0.inst_src_2_ ),
    .C(execution_unit_0.gie ),
    .Y(_03086_)
  );
  NAND2X1 _08532_ (
    .A(execution_unit_0.register_file_0.r12_3_ ),
    .B(_03011_),
    .Y(_03087_)
  );
  NAND2X1 _08533_ (
    .A(execution_unit_0.register_file_0.r5_3_ ),
    .B(_03004_),
    .Y(_03088_)
  );
  AOI22X1 _08534_ (
    .A(execution_unit_0.register_file_0.r11_3_ ),
    .B(_03009_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_3_ ),
    .Y(_03089_)
  );
  AOI22X1 _08535_ (
    .A(execution_unit_0.register_file_0.r14_3_ ),
    .B(_02997_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_3_ ),
    .Y(_03090_)
  );
  NAND3X1 _08536_ (
    .A(_03087_),
    .B(_03089_),
    .C(_03090_),
    .Y(_03091_)
  );
  AOI22X1 _08537_ (
    .A(execution_unit_0.register_file_0.r1_3_ ),
    .B(_03001_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_3_ ),
    .Y(_03092_)
  );
  AOI22X1 _08538_ (
    .A(dbg_0.UNUSED_pc_3_ ),
    .B(_03015_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_3_ ),
    .Y(_03093_)
  );
  NAND3X1 _08539_ (
    .A(_03088_),
    .B(_03092_),
    .C(_03093_),
    .Y(_03094_)
  );
  NOR2X1 _08540_ (
    .A(_03091_),
    .B(_03094_),
    .Y(_03095_)
  );
  AOI22X1 _08541_ (
    .A(execution_unit_0.register_file_0.r13_3_ ),
    .B(_02990_),
    .C(_02995_),
    .D(execution_unit_0.register_file_0.r7_3_ ),
    .Y(_03096_)
  );
  OAI21X1 _08542_ (
    .A(_02960_),
    .B(_02993_),
    .C(_03096_),
    .Y(_03097_)
  );
  AOI22X1 _08543_ (
    .A(execution_unit_0.register_file_0.r3_3_ ),
    .B(_03005_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_3_ ),
    .Y(_03098_)
  );
  NAND2X1 _08544_ (
    .A(_03086_),
    .B(_03098_),
    .Y(_03099_)
  );
  NOR2X1 _08545_ (
    .A(_03097_),
    .B(_03099_),
    .Y(_03100_)
  );
  AND2X1 _08546_ (
    .A(_03095_),
    .B(_03100_),
    .Y(_03101_)
  );
  INVX1 _08547_ (
    .A(_03101_),
    .Y(execution_unit_0.reg_src_3_ )
  );
  NOR3X1 _08548_ (
    .A(_03061_),
    .B(_03081_),
    .C(_03101_),
    .Y(_03102_)
  );
  NOR2X1 _08549_ (
    .A(_03082_),
    .B(execution_unit_0.reg_src_3_ ),
    .Y(_03103_)
  );
  NOR2X1 _08550_ (
    .A(_03102_),
    .B(_03103_),
    .Y(_03104_)
  );
  NOR2X1 _08551_ (
    .A(execution_unit_0.register_file_0.r15_3_ ),
    .B(_03033_),
    .Y(_03105_)
  );
  OAI21X1 _08552_ (
    .A(_03034_),
    .B(_03104_),
    .C(_03032_),
    .Y(_03106_)
  );
  OAI22X1 _08553_ (
    .A(_02962_),
    .B(_03032_),
    .C(_03105_),
    .D(_03106_),
    .Y(_02009_)
  );
  AOI22X1 _08554_ (
    .A(execution_unit_0.register_file_0.r10_4_ ),
    .B(_02992_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_4_ ),
    .Y(_03107_)
  );
  AOI22X1 _08555_ (
    .A(dbg_0.UNUSED_pc_4_ ),
    .B(_03015_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_4_ ),
    .Y(_03108_)
  );
  NAND2X1 _08556_ (
    .A(_03107_),
    .B(_03108_),
    .Y(_03109_)
  );
  AOI22X1 _08557_ (
    .A(execution_unit_0.register_file_0.r11_4_ ),
    .B(_03009_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_4_ ),
    .Y(_03110_)
  );
  AOI22X1 _08558_ (
    .A(execution_unit_0.register_file_0.r3_4_ ),
    .B(_03005_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_4_ ),
    .Y(_03111_)
  );
  NAND2X1 _08559_ (
    .A(_03110_),
    .B(_03111_),
    .Y(_03112_)
  );
  NOR2X1 _08560_ (
    .A(_03109_),
    .B(_03112_),
    .Y(_03113_)
  );
  AOI22X1 _08561_ (
    .A(execution_unit_0.register_file_0.r1_4_ ),
    .B(_03001_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_4_ ),
    .Y(_03114_)
  );
  AOI22X1 _08562_ (
    .A(execution_unit_0.register_file_0.r7_4_ ),
    .B(_02995_),
    .C(_03004_),
    .D(execution_unit_0.register_file_0.r5_4_ ),
    .Y(_03115_)
  );
  NAND2X1 _08563_ (
    .A(_03114_),
    .B(_03115_),
    .Y(_03116_)
  );
  AOI22X1 _08564_ (
    .A(execution_unit_0.register_file_0.r14_4_ ),
    .B(_02997_),
    .C(_02999_),
    .D(execution_unit_0.register_file_0.r2_4_ ),
    .Y(_03117_)
  );
  AOI22X1 _08565_ (
    .A(execution_unit_0.register_file_0.r13_4_ ),
    .B(_02990_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_4_ ),
    .Y(_03118_)
  );
  NAND2X1 _08566_ (
    .A(_03117_),
    .B(_03118_),
    .Y(_03119_)
  );
  NOR2X1 _08567_ (
    .A(_03116_),
    .B(_03119_),
    .Y(_03120_)
  );
  NAND2X1 _08568_ (
    .A(_03113_),
    .B(_03120_),
    .Y(execution_unit_0.reg_src_4_ )
  );
  NAND2X1 _08569_ (
    .A(_03102_),
    .B(execution_unit_0.reg_src_4_ ),
    .Y(_03121_)
  );
  XOR2X1 _08570_ (
    .A(_03102_),
    .B(execution_unit_0.reg_src_4_ ),
    .Y(_03122_)
  );
  NOR2X1 _08571_ (
    .A(execution_unit_0.register_file_0.r15_4_ ),
    .B(_03033_),
    .Y(_03123_)
  );
  OAI21X1 _08572_ (
    .A(_03034_),
    .B(_03122_),
    .C(_03032_),
    .Y(_03124_)
  );
  OAI22X1 _08573_ (
    .A(_02965_),
    .B(_03032_),
    .C(_03123_),
    .D(_03124_),
    .Y(_02010_)
  );
  AOI22X1 _08574_ (
    .A(execution_unit_0.register_file_0.r7_5_ ),
    .B(_02995_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_5_ ),
    .Y(_03125_)
  );
  AOI22X1 _08575_ (
    .A(execution_unit_0.register_file_0.r3_5_ ),
    .B(_03005_),
    .C(_03009_),
    .D(execution_unit_0.register_file_0.r11_5_ ),
    .Y(_03126_)
  );
  NAND2X1 _08576_ (
    .A(_03125_),
    .B(_03126_),
    .Y(_03127_)
  );
  AOI22X1 _08577_ (
    .A(execution_unit_0.register_file_0.r13_5_ ),
    .B(_02990_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_5_ ),
    .Y(_03128_)
  );
  AOI22X1 _08578_ (
    .A(execution_unit_0.register_file_0.r10_5_ ),
    .B(_02992_),
    .C(_02997_),
    .D(execution_unit_0.register_file_0.r14_5_ ),
    .Y(_03129_)
  );
  NAND2X1 _08579_ (
    .A(_03128_),
    .B(_03129_),
    .Y(_03130_)
  );
  NOR2X1 _08580_ (
    .A(_03127_),
    .B(_03130_),
    .Y(_03131_)
  );
  AOI22X1 _08581_ (
    .A(execution_unit_0.register_file_0.r12_5_ ),
    .B(_03011_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_5_ ),
    .Y(_03132_)
  );
  AOI22X1 _08582_ (
    .A(execution_unit_0.register_file_0.r5_5_ ),
    .B(_03004_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_5_ ),
    .Y(_03133_)
  );
  NAND2X1 _08583_ (
    .A(_03132_),
    .B(_03133_),
    .Y(_03134_)
  );
  AOI22X1 _08584_ (
    .A(execution_unit_0.register_file_0.r1_5_ ),
    .B(_03001_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_5_ ),
    .Y(_03135_)
  );
  AOI22X1 _08585_ (
    .A(clock_module_0.oscoff ),
    .B(_02999_),
    .C(_03015_),
    .D(dbg_0.UNUSED_pc_5_ ),
    .Y(_03136_)
  );
  NAND2X1 _08586_ (
    .A(_03135_),
    .B(_03136_),
    .Y(_03137_)
  );
  NOR2X1 _08587_ (
    .A(_03134_),
    .B(_03137_),
    .Y(_03138_)
  );
  NAND2X1 _08588_ (
    .A(_03131_),
    .B(_03138_),
    .Y(execution_unit_0.reg_src_5_ )
  );
  NAND3X1 _08589_ (
    .A(_03102_),
    .B(execution_unit_0.reg_src_4_ ),
    .C(execution_unit_0.reg_src_5_ ),
    .Y(_03139_)
  );
  XNOR2X1 _08590_ (
    .A(_03121_),
    .B(execution_unit_0.reg_src_5_ ),
    .Y(_03140_)
  );
  NOR2X1 _08591_ (
    .A(execution_unit_0.register_file_0.r15_5_ ),
    .B(_03033_),
    .Y(_03141_)
  );
  OAI21X1 _08592_ (
    .A(_03034_),
    .B(_03140_),
    .C(_03032_),
    .Y(_03142_)
  );
  OAI22X1 _08593_ (
    .A(_02966_),
    .B(_03032_),
    .C(_03141_),
    .D(_03142_),
    .Y(_02011_)
  );
  AOI22X1 _08594_ (
    .A(execution_unit_0.register_file_0.r5_6_ ),
    .B(_03004_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_6_ ),
    .Y(_03143_)
  );
  AOI22X1 _08595_ (
    .A(execution_unit_0.register_file_0.r14_6_ ),
    .B(_02997_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_6_ ),
    .Y(_03144_)
  );
  AND2X1 _08596_ (
    .A(_03143_),
    .B(_03144_),
    .Y(_03145_)
  );
  AOI22X1 _08597_ (
    .A(execution_unit_0.register_file_0.r3_6_ ),
    .B(_03005_),
    .C(_03009_),
    .D(execution_unit_0.register_file_0.r11_6_ ),
    .Y(_03146_)
  );
  AOI22X1 _08598_ (
    .A(execution_unit_0.register_file_0.r7_6_ ),
    .B(_02995_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_6_ ),
    .Y(_03147_)
  );
  NAND3X1 _08599_ (
    .A(_03145_),
    .B(_03146_),
    .C(_03147_),
    .Y(_03148_)
  );
  AOI22X1 _08600_ (
    .A(execution_unit_0.register_file_0.r10_6_ ),
    .B(_02992_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_6_ ),
    .Y(_03149_)
  );
  INVX1 _08601_ (
    .A(_03149_),
    .Y(_03150_)
  );
  AOI21X1 _08602_ (
    .A(execution_unit_0.register_file_0.r1_6_ ),
    .B(_03001_),
    .C(_03150_),
    .Y(_03151_)
  );
  AOI22X1 _08603_ (
    .A(execution_unit_0.register_file_0.r13_6_ ),
    .B(_02990_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_6_ ),
    .Y(_03152_)
  );
  AOI22X1 _08604_ (
    .A(execution_unit_0.register_file_0.r6_6_ ),
    .B(_03013_),
    .C(_03015_),
    .D(dbg_0.UNUSED_pc_6_ ),
    .Y(_03153_)
  );
  NAND3X1 _08605_ (
    .A(_03151_),
    .B(_03152_),
    .C(_03153_),
    .Y(_03154_)
  );
  OR2X1 _08606_ (
    .A(_03148_),
    .B(_03154_),
    .Y(execution_unit_0.reg_src_6_ )
  );
  INVX1 _08607_ (
    .A(execution_unit_0.reg_src_6_ ),
    .Y(_03155_)
  );
  NOR2X1 _08608_ (
    .A(_03139_),
    .B(_03155_),
    .Y(_03156_)
  );
  XNOR2X1 _08609_ (
    .A(_03139_),
    .B(_03155_),
    .Y(_03157_)
  );
  AOI21X1 _08610_ (
    .A(_03033_),
    .B(_03157_),
    .C(_03031_),
    .Y(_03158_)
  );
  OAI21X1 _08611_ (
    .A(execution_unit_0.register_file_0.r15_6_ ),
    .B(_03033_),
    .C(_03158_),
    .Y(_03159_)
  );
  OAI21X1 _08612_ (
    .A(_02967_),
    .B(_03032_),
    .C(_03159_),
    .Y(_02012_)
  );
  AOI22X1 _08613_ (
    .A(dbg_0.UNUSED_pc_7_ ),
    .B(_03015_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_7_ ),
    .Y(_03160_)
  );
  AOI22X1 _08614_ (
    .A(execution_unit_0.register_file_0.r5_7_ ),
    .B(_03004_),
    .C(_03005_),
    .D(execution_unit_0.register_file_0.r3_7_ ),
    .Y(_03161_)
  );
  NAND2X1 _08615_ (
    .A(_03160_),
    .B(_03161_),
    .Y(_03162_)
  );
  AOI22X1 _08616_ (
    .A(execution_unit_0.register_file_0.r14_7_ ),
    .B(_02997_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_7_ ),
    .Y(_03163_)
  );
  AOI22X1 _08617_ (
    .A(execution_unit_0.register_file_0.r13_7_ ),
    .B(_02990_),
    .C(_02992_),
    .D(execution_unit_0.register_file_0.r10_7_ ),
    .Y(_03164_)
  );
  NAND2X1 _08618_ (
    .A(_03163_),
    .B(_03164_),
    .Y(_03165_)
  );
  NOR2X1 _08619_ (
    .A(_03162_),
    .B(_03165_),
    .Y(_03166_)
  );
  AOI22X1 _08620_ (
    .A(execution_unit_0.register_file_0.r1_7_ ),
    .B(_03001_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_7_ ),
    .Y(_03167_)
  );
  AOI22X1 _08621_ (
    .A(clock_module_0.scg1 ),
    .B(_02999_),
    .C(_03009_),
    .D(execution_unit_0.register_file_0.r11_7_ ),
    .Y(_03168_)
  );
  NAND2X1 _08622_ (
    .A(_03167_),
    .B(_03168_),
    .Y(_03169_)
  );
  AOI22X1 _08623_ (
    .A(execution_unit_0.register_file_0.r7_7_ ),
    .B(_02995_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_7_ ),
    .Y(_03170_)
  );
  AOI22X1 _08624_ (
    .A(execution_unit_0.register_file_0.r6_7_ ),
    .B(_03013_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_7_ ),
    .Y(_03171_)
  );
  NAND2X1 _08625_ (
    .A(_03170_),
    .B(_03171_),
    .Y(_03172_)
  );
  NOR2X1 _08626_ (
    .A(_03169_),
    .B(_03172_),
    .Y(_03173_)
  );
  NAND2X1 _08627_ (
    .A(_03166_),
    .B(_03173_),
    .Y(execution_unit_0.reg_src_7_ )
  );
  INVX1 _08628_ (
    .A(execution_unit_0.reg_src_7_ ),
    .Y(_03174_)
  );
  NOR3X1 _08629_ (
    .A(_03139_),
    .B(_03155_),
    .C(_03174_),
    .Y(_03175_)
  );
  NOR2X1 _08630_ (
    .A(_03156_),
    .B(execution_unit_0.reg_src_7_ ),
    .Y(_03176_)
  );
  NOR2X1 _08631_ (
    .A(_03175_),
    .B(_03176_),
    .Y(_03177_)
  );
  NOR2X1 _08632_ (
    .A(execution_unit_0.register_file_0.r15_7_ ),
    .B(_03033_),
    .Y(_03178_)
  );
  OAI21X1 _08633_ (
    .A(_03034_),
    .B(_03177_),
    .C(_03032_),
    .Y(_03179_)
  );
  OAI22X1 _08634_ (
    .A(_02968_),
    .B(_03032_),
    .C(_03178_),
    .D(_03179_),
    .Y(_02013_)
  );
  NAND2X1 _08635_ (
    .A(execution_unit_0.register_file_0.r14_8_ ),
    .B(_02997_),
    .Y(_03180_)
  );
  OAI21X1 _08636_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(execution_unit_0.inst_src_2_ ),
    .C(execution_unit_0.alu_0.status_3_ ),
    .Y(_03181_)
  );
  AOI22X1 _08637_ (
    .A(execution_unit_0.register_file_0.r4_8_ ),
    .B(_03007_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_8_ ),
    .Y(_03182_)
  );
  AOI22X1 _08638_ (
    .A(execution_unit_0.register_file_0.r5_8_ ),
    .B(_03004_),
    .C(_03015_),
    .D(dbg_0.UNUSED_pc_8_ ),
    .Y(_03183_)
  );
  AOI22X1 _08639_ (
    .A(execution_unit_0.register_file_0.r13_8_ ),
    .B(_02990_),
    .C(_02995_),
    .D(execution_unit_0.register_file_0.r7_8_ ),
    .Y(_03184_)
  );
  NAND2X1 _08640_ (
    .A(_03180_),
    .B(_03184_),
    .Y(_03185_)
  );
  AOI21X1 _08641_ (
    .A(execution_unit_0.register_file_0.r11_8_ ),
    .B(_03009_),
    .C(_03185_),
    .Y(_03186_)
  );
  NAND3X1 _08642_ (
    .A(_03182_),
    .B(_03183_),
    .C(_03186_),
    .Y(_03187_)
  );
  AOI22X1 _08643_ (
    .A(execution_unit_0.register_file_0.r3_8_ ),
    .B(_03005_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_8_ ),
    .Y(_03188_)
  );
  AOI22X1 _08644_ (
    .A(execution_unit_0.register_file_0.r1_8_ ),
    .B(_03001_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_8_ ),
    .Y(_03189_)
  );
  AOI22X1 _08645_ (
    .A(execution_unit_0.register_file_0.r10_8_ ),
    .B(_02992_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_8_ ),
    .Y(_03190_)
  );
  NAND2X1 _08646_ (
    .A(_03189_),
    .B(_03190_),
    .Y(_03191_)
  );
  AOI21X1 _08647_ (
    .A(execution_unit_0.register_file_0.r8_8_ ),
    .B(_03022_),
    .C(_03191_),
    .Y(_03192_)
  );
  NAND3X1 _08648_ (
    .A(_03181_),
    .B(_03188_),
    .C(_03192_),
    .Y(_03193_)
  );
  OR2X1 _08649_ (
    .A(_03187_),
    .B(_03193_),
    .Y(execution_unit_0.reg_src_8_ )
  );
  OAI21X1 _08650_ (
    .A(_03187_),
    .B(_03193_),
    .C(_03175_),
    .Y(_03194_)
  );
  XOR2X1 _08651_ (
    .A(_03175_),
    .B(execution_unit_0.reg_src_8_ ),
    .Y(_03195_)
  );
  OAI21X1 _08652_ (
    .A(_03034_),
    .B(_03195_),
    .C(_03032_),
    .Y(_03196_)
  );
  INVX1 _08653_ (
    .A(_03196_),
    .Y(_03197_)
  );
  OAI21X1 _08654_ (
    .A(execution_unit_0.register_file_0.r15_8_ ),
    .B(_03033_),
    .C(_03197_),
    .Y(_03198_)
  );
  OAI21X1 _08655_ (
    .A(_02982_),
    .B(_03032_),
    .C(_03198_),
    .Y(_02014_)
  );
  AOI22X1 _08656_ (
    .A(execution_unit_0.register_file_0.r10_9_ ),
    .B(_02992_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_9_ ),
    .Y(_03199_)
  );
  AOI22X1 _08657_ (
    .A(execution_unit_0.register_file_0.r14_9_ ),
    .B(_02997_),
    .C(_03001_),
    .D(execution_unit_0.register_file_0.r1_9_ ),
    .Y(_03200_)
  );
  AND2X1 _08658_ (
    .A(_03199_),
    .B(_03200_),
    .Y(_03201_)
  );
  AOI22X1 _08659_ (
    .A(execution_unit_0.register_file_0.r7_9_ ),
    .B(_02995_),
    .C(_03004_),
    .D(execution_unit_0.register_file_0.r5_9_ ),
    .Y(_03202_)
  );
  AOI22X1 _08660_ (
    .A(execution_unit_0.register_file_0.r3_9_ ),
    .B(_03005_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_9_ ),
    .Y(_03203_)
  );
  NAND3X1 _08661_ (
    .A(_03201_),
    .B(_03202_),
    .C(_03203_),
    .Y(_03204_)
  );
  AOI22X1 _08662_ (
    .A(execution_unit_0.register_file_0.r11_9_ ),
    .B(_03009_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_9_ ),
    .Y(_03205_)
  );
  INVX1 _08663_ (
    .A(_03205_),
    .Y(_03206_)
  );
  AOI21X1 _08664_ (
    .A(execution_unit_0.register_file_0.r8_9_ ),
    .B(_03022_),
    .C(_03206_),
    .Y(_03207_)
  );
  AOI22X1 _08665_ (
    .A(execution_unit_0.register_file_0.r12_9_ ),
    .B(_03011_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_9_ ),
    .Y(_03208_)
  );
  AOI22X1 _08666_ (
    .A(execution_unit_0.register_file_0.r13_9_ ),
    .B(_02990_),
    .C(_03015_),
    .D(dbg_0.UNUSED_pc_9_ ),
    .Y(_03209_)
  );
  NAND3X1 _08667_ (
    .A(_03207_),
    .B(_03208_),
    .C(_03209_),
    .Y(_03210_)
  );
  OR2X1 _08668_ (
    .A(_03204_),
    .B(_03210_),
    .Y(execution_unit_0.reg_src_9_ )
  );
  NAND3X1 _08669_ (
    .A(_03175_),
    .B(execution_unit_0.reg_src_8_ ),
    .C(execution_unit_0.reg_src_9_ ),
    .Y(_03211_)
  );
  XNOR2X1 _08670_ (
    .A(_03194_),
    .B(execution_unit_0.reg_src_9_ ),
    .Y(_03212_)
  );
  OAI21X1 _08671_ (
    .A(_03034_),
    .B(_03212_),
    .C(_03032_),
    .Y(_03213_)
  );
  INVX1 _08672_ (
    .A(_03213_),
    .Y(_03214_)
  );
  OAI21X1 _08673_ (
    .A(execution_unit_0.register_file_0.r15_9_ ),
    .B(_03033_),
    .C(_03214_),
    .Y(_03215_)
  );
  OAI21X1 _08674_ (
    .A(_02983_),
    .B(_03032_),
    .C(_03215_),
    .Y(_02015_)
  );
  NAND2X1 _08675_ (
    .A(execution_unit_0.register_file_0.r9_10_ ),
    .B(_03017_),
    .Y(_03216_)
  );
  NAND2X1 _08676_ (
    .A(execution_unit_0.register_file_0.r7_10_ ),
    .B(_02995_),
    .Y(_03217_)
  );
  AOI22X1 _08677_ (
    .A(execution_unit_0.register_file_0.r5_10_ ),
    .B(_03004_),
    .C(_03015_),
    .D(dbg_0.UNUSED_pc_10_ ),
    .Y(_03218_)
  );
  NAND2X1 _08678_ (
    .A(_03217_),
    .B(_03218_),
    .Y(_03219_)
  );
  AOI22X1 _08679_ (
    .A(execution_unit_0.register_file_0.r4_10_ ),
    .B(_03007_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_10_ ),
    .Y(_03220_)
  );
  AOI22X1 _08680_ (
    .A(execution_unit_0.register_file_0.r13_10_ ),
    .B(_02990_),
    .C(_03001_),
    .D(execution_unit_0.register_file_0.r1_10_ ),
    .Y(_03221_)
  );
  NAND3X1 _08681_ (
    .A(_03216_),
    .B(_03220_),
    .C(_03221_),
    .Y(_03222_)
  );
  NOR2X1 _08682_ (
    .A(_03219_),
    .B(_03222_),
    .Y(_03223_)
  );
  AOI22X1 _08683_ (
    .A(execution_unit_0.register_file_0.r11_10_ ),
    .B(_03009_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_10_ ),
    .Y(_03224_)
  );
  AOI22X1 _08684_ (
    .A(execution_unit_0.register_file_0.r10_10_ ),
    .B(_02992_),
    .C(_03005_),
    .D(execution_unit_0.register_file_0.r3_10_ ),
    .Y(_03225_)
  );
  AOI22X1 _08685_ (
    .A(execution_unit_0.register_file_0.r14_10_ ),
    .B(_02997_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_10_ ),
    .Y(_03226_)
  );
  NAND3X1 _08686_ (
    .A(_03224_),
    .B(_03225_),
    .C(_03226_),
    .Y(_03227_)
  );
  AOI21X1 _08687_ (
    .A(execution_unit_0.register_file_0.r8_10_ ),
    .B(_03022_),
    .C(_03227_),
    .Y(_03228_)
  );
  NAND2X1 _08688_ (
    .A(_03223_),
    .B(_03228_),
    .Y(execution_unit_0.reg_src_10_ )
  );
  INVX1 _08689_ (
    .A(execution_unit_0.reg_src_10_ ),
    .Y(_03229_)
  );
  NOR2X1 _08690_ (
    .A(_03211_),
    .B(_03229_),
    .Y(_03230_)
  );
  XNOR2X1 _08691_ (
    .A(_03211_),
    .B(_03229_),
    .Y(_03231_)
  );
  AOI21X1 _08692_ (
    .A(_03033_),
    .B(_03231_),
    .C(_03031_),
    .Y(_03232_)
  );
  OAI21X1 _08693_ (
    .A(execution_unit_0.register_file_0.r15_10_ ),
    .B(_03033_),
    .C(_03232_),
    .Y(_03233_)
  );
  OAI21X1 _08694_ (
    .A(_02984_),
    .B(_03032_),
    .C(_03233_),
    .Y(_02001_)
  );
  AOI22X1 _08695_ (
    .A(execution_unit_0.register_file_0.r14_11_ ),
    .B(_02997_),
    .C(_03001_),
    .D(execution_unit_0.register_file_0.r1_11_ ),
    .Y(_03234_)
  );
  AOI22X1 _08696_ (
    .A(execution_unit_0.register_file_0.r9_11_ ),
    .B(_03017_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_11_ ),
    .Y(_03235_)
  );
  AND2X1 _08697_ (
    .A(_03234_),
    .B(_03235_),
    .Y(_03236_)
  );
  AOI22X1 _08698_ (
    .A(execution_unit_0.register_file_0.r10_11_ ),
    .B(_02992_),
    .C(_02995_),
    .D(execution_unit_0.register_file_0.r7_11_ ),
    .Y(_03237_)
  );
  AOI22X1 _08699_ (
    .A(execution_unit_0.register_file_0.r13_11_ ),
    .B(_02990_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_11_ ),
    .Y(_03238_)
  );
  NAND3X1 _08700_ (
    .A(_03236_),
    .B(_03237_),
    .C(_03238_),
    .Y(_03239_)
  );
  AOI22X1 _08701_ (
    .A(execution_unit_0.register_file_0.r5_11_ ),
    .B(_03004_),
    .C(_03009_),
    .D(execution_unit_0.register_file_0.r11_11_ ),
    .Y(_03240_)
  );
  INVX1 _08702_ (
    .A(_03240_),
    .Y(_03241_)
  );
  AOI21X1 _08703_ (
    .A(dbg_0.UNUSED_pc_11_ ),
    .B(_03015_),
    .C(_03241_),
    .Y(_03242_)
  );
  AOI22X1 _08704_ (
    .A(execution_unit_0.register_file_0.r3_11_ ),
    .B(_03005_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_11_ ),
    .Y(_03243_)
  );
  AOI22X1 _08705_ (
    .A(execution_unit_0.register_file_0.r4_11_ ),
    .B(_03007_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_11_ ),
    .Y(_03244_)
  );
  NAND3X1 _08706_ (
    .A(_03242_),
    .B(_03243_),
    .C(_03244_),
    .Y(_03245_)
  );
  OR2X1 _08707_ (
    .A(_03239_),
    .B(_03245_),
    .Y(execution_unit_0.reg_src_11_ )
  );
  INVX1 _08708_ (
    .A(execution_unit_0.reg_src_11_ ),
    .Y(_03246_)
  );
  NOR3X1 _08709_ (
    .A(_03211_),
    .B(_03229_),
    .C(_03246_),
    .Y(_03247_)
  );
  NOR2X1 _08710_ (
    .A(_03230_),
    .B(execution_unit_0.reg_src_11_ ),
    .Y(_03248_)
  );
  NOR2X1 _08711_ (
    .A(_03247_),
    .B(_03248_),
    .Y(_03249_)
  );
  OAI21X1 _08712_ (
    .A(execution_unit_0.register_file_0.r15_11_ ),
    .B(_03033_),
    .C(_03032_),
    .Y(_03250_)
  );
  INVX1 _08713_ (
    .A(_03250_),
    .Y(_03251_)
  );
  OAI21X1 _08714_ (
    .A(_03034_),
    .B(_03249_),
    .C(_03251_),
    .Y(_03252_)
  );
  OAI21X1 _08715_ (
    .A(_02985_),
    .B(_03032_),
    .C(_03252_),
    .Y(_02002_)
  );
  NAND2X1 _08716_ (
    .A(dbg_0.UNUSED_pc_12_ ),
    .B(_03015_),
    .Y(_03253_)
  );
  AOI22X1 _08717_ (
    .A(execution_unit_0.register_file_0.r14_12_ ),
    .B(_02997_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_12_ ),
    .Y(_03254_)
  );
  NAND2X1 _08718_ (
    .A(execution_unit_0.register_file_0.r5_12_ ),
    .B(_03004_),
    .Y(_03255_)
  );
  AOI22X1 _08719_ (
    .A(execution_unit_0.register_file_0.r3_12_ ),
    .B(_03005_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_12_ ),
    .Y(_03256_)
  );
  AOI22X1 _08720_ (
    .A(execution_unit_0.register_file_0.r6_12_ ),
    .B(_03013_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_12_ ),
    .Y(_03257_)
  );
  AOI22X1 _08721_ (
    .A(execution_unit_0.register_file_0.r10_12_ ),
    .B(_02992_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_12_ ),
    .Y(_03258_)
  );
  NAND3X1 _08722_ (
    .A(_03256_),
    .B(_03257_),
    .C(_03258_),
    .Y(_03259_)
  );
  AOI21X1 _08723_ (
    .A(execution_unit_0.register_file_0.r11_12_ ),
    .B(_03009_),
    .C(_03259_),
    .Y(_03260_)
  );
  AOI22X1 _08724_ (
    .A(execution_unit_0.register_file_0.r13_12_ ),
    .B(_02990_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_12_ ),
    .Y(_03261_)
  );
  NAND2X1 _08725_ (
    .A(_03253_),
    .B(_03261_),
    .Y(_03262_)
  );
  AOI22X1 _08726_ (
    .A(execution_unit_0.register_file_0.r7_12_ ),
    .B(_02995_),
    .C(_03001_),
    .D(execution_unit_0.register_file_0.r1_12_ ),
    .Y(_03263_)
  );
  NAND2X1 _08727_ (
    .A(_03255_),
    .B(_03263_),
    .Y(_03264_)
  );
  NOR2X1 _08728_ (
    .A(_03262_),
    .B(_03264_),
    .Y(_03265_)
  );
  NAND3X1 _08729_ (
    .A(_03254_),
    .B(_03260_),
    .C(_03265_),
    .Y(execution_unit_0.reg_src_12_ )
  );
  NAND2X1 _08730_ (
    .A(_03247_),
    .B(execution_unit_0.reg_src_12_ ),
    .Y(_03266_)
  );
  XOR2X1 _08731_ (
    .A(_03247_),
    .B(execution_unit_0.reg_src_12_ ),
    .Y(_03267_)
  );
  OAI21X1 _08732_ (
    .A(execution_unit_0.register_file_0.r15_12_ ),
    .B(_03033_),
    .C(_03032_),
    .Y(_03268_)
  );
  INVX1 _08733_ (
    .A(_03268_),
    .Y(_03269_)
  );
  OAI21X1 _08734_ (
    .A(_03034_),
    .B(_03267_),
    .C(_03269_),
    .Y(_03270_)
  );
  OAI21X1 _08735_ (
    .A(_02986_),
    .B(_03032_),
    .C(_03270_),
    .Y(_02003_)
  );
  NAND2X1 _08736_ (
    .A(execution_unit_0.register_file_0.r5_13_ ),
    .B(_03004_),
    .Y(_03271_)
  );
  AOI22X1 _08737_ (
    .A(execution_unit_0.register_file_0.r15_13_ ),
    .B(_03020_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_13_ ),
    .Y(_03272_)
  );
  NAND2X1 _08738_ (
    .A(_03271_),
    .B(_03272_),
    .Y(_03273_)
  );
  AOI21X1 _08739_ (
    .A(execution_unit_0.register_file_0.r14_13_ ),
    .B(_02997_),
    .C(_03273_),
    .Y(_03274_)
  );
  AOI22X1 _08740_ (
    .A(execution_unit_0.register_file_0.r13_13_ ),
    .B(_02990_),
    .C(_03001_),
    .D(execution_unit_0.register_file_0.r1_13_ ),
    .Y(_03275_)
  );
  AOI22X1 _08741_ (
    .A(execution_unit_0.register_file_0.r3_13_ ),
    .B(_03005_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_13_ ),
    .Y(_03276_)
  );
  NAND3X1 _08742_ (
    .A(_03274_),
    .B(_03275_),
    .C(_03276_),
    .Y(_03277_)
  );
  INVX1 _08743_ (
    .A(_03277_),
    .Y(_03278_)
  );
  AOI22X1 _08744_ (
    .A(execution_unit_0.register_file_0.r11_13_ ),
    .B(_03009_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_13_ ),
    .Y(_03279_)
  );
  AOI22X1 _08745_ (
    .A(execution_unit_0.register_file_0.r7_13_ ),
    .B(_02995_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_13_ ),
    .Y(_03280_)
  );
  AOI22X1 _08746_ (
    .A(execution_unit_0.register_file_0.r10_13_ ),
    .B(_02992_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_13_ ),
    .Y(_03281_)
  );
  NAND2X1 _08747_ (
    .A(_03280_),
    .B(_03281_),
    .Y(_03282_)
  );
  AOI21X1 _08748_ (
    .A(dbg_0.UNUSED_pc_13_ ),
    .B(_03015_),
    .C(_03282_),
    .Y(_03283_)
  );
  NAND3X1 _08749_ (
    .A(_03278_),
    .B(_03279_),
    .C(_03283_),
    .Y(execution_unit_0.reg_src_13_ )
  );
  NAND3X1 _08750_ (
    .A(_03247_),
    .B(execution_unit_0.reg_src_12_ ),
    .C(execution_unit_0.reg_src_13_ ),
    .Y(_03284_)
  );
  XNOR2X1 _08751_ (
    .A(_03266_),
    .B(execution_unit_0.reg_src_13_ ),
    .Y(_03285_)
  );
  OAI21X1 _08752_ (
    .A(execution_unit_0.register_file_0.r15_13_ ),
    .B(_03033_),
    .C(_03032_),
    .Y(_03286_)
  );
  INVX1 _08753_ (
    .A(_03286_),
    .Y(_03287_)
  );
  OAI21X1 _08754_ (
    .A(_03034_),
    .B(_03285_),
    .C(_03287_),
    .Y(_03288_)
  );
  OAI21X1 _08755_ (
    .A(_02987_),
    .B(_03032_),
    .C(_03288_),
    .Y(_02004_)
  );
  NAND2X1 _08756_ (
    .A(execution_unit_0.register_file_0.r8_14_ ),
    .B(_03022_),
    .Y(_03289_)
  );
  AOI22X1 _08757_ (
    .A(execution_unit_0.register_file_0.r10_14_ ),
    .B(_02992_),
    .C(_03009_),
    .D(execution_unit_0.register_file_0.r11_14_ ),
    .Y(_03290_)
  );
  AOI22X1 _08758_ (
    .A(execution_unit_0.register_file_0.r14_14_ ),
    .B(_02997_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_14_ ),
    .Y(_03291_)
  );
  AOI22X1 _08759_ (
    .A(execution_unit_0.register_file_0.r13_14_ ),
    .B(_02990_),
    .C(_03020_),
    .D(execution_unit_0.register_file_0.r15_14_ ),
    .Y(_03292_)
  );
  NAND3X1 _08760_ (
    .A(_03290_),
    .B(_03291_),
    .C(_03292_),
    .Y(_03293_)
  );
  AOI21X1 _08761_ (
    .A(execution_unit_0.register_file_0.r1_14_ ),
    .B(_03001_),
    .C(_03293_),
    .Y(_03294_)
  );
  AOI22X1 _08762_ (
    .A(execution_unit_0.register_file_0.r7_14_ ),
    .B(_02995_),
    .C(_03015_),
    .D(dbg_0.UNUSED_pc_14_ ),
    .Y(_03295_)
  );
  AOI22X1 _08763_ (
    .A(execution_unit_0.register_file_0.r5_14_ ),
    .B(_03004_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_14_ ),
    .Y(_03296_)
  );
  NAND2X1 _08764_ (
    .A(_03289_),
    .B(_03296_),
    .Y(_03297_)
  );
  AOI22X1 _08765_ (
    .A(execution_unit_0.register_file_0.r3_14_ ),
    .B(_03005_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_14_ ),
    .Y(_03298_)
  );
  OAI21X1 _08766_ (
    .A(_02972_),
    .B(_03018_),
    .C(_03298_),
    .Y(_03299_)
  );
  NOR2X1 _08767_ (
    .A(_03297_),
    .B(_03299_),
    .Y(_03300_)
  );
  NAND3X1 _08768_ (
    .A(_03294_),
    .B(_03295_),
    .C(_03300_),
    .Y(execution_unit_0.reg_src_14_ )
  );
  INVX1 _08769_ (
    .A(execution_unit_0.reg_src_14_ ),
    .Y(_03301_)
  );
  NOR2X1 _08770_ (
    .A(_03284_),
    .B(_03301_),
    .Y(_03302_)
  );
  XNOR2X1 _08771_ (
    .A(_03284_),
    .B(execution_unit_0.reg_src_14_ ),
    .Y(_03303_)
  );
  OAI21X1 _08772_ (
    .A(execution_unit_0.register_file_0.r15_14_ ),
    .B(_03033_),
    .C(_03032_),
    .Y(_03304_)
  );
  INVX1 _08773_ (
    .A(_03304_),
    .Y(_03305_)
  );
  OAI21X1 _08774_ (
    .A(_03034_),
    .B(_03303_),
    .C(_03305_),
    .Y(_03306_)
  );
  OAI21X1 _08775_ (
    .A(_02988_),
    .B(_03032_),
    .C(_03306_),
    .Y(_02005_)
  );
  AOI22X1 _08776_ (
    .A(execution_unit_0.register_file_0.r11_15_ ),
    .B(_03009_),
    .C(_03013_),
    .D(execution_unit_0.register_file_0.r6_15_ ),
    .Y(_02153_)
  );
  NAND2X1 _08777_ (
    .A(execution_unit_0.register_file_0.r1_15_ ),
    .B(_03001_),
    .Y(_02154_)
  );
  AOI22X1 _08778_ (
    .A(execution_unit_0.register_file_0.r5_15_ ),
    .B(_03004_),
    .C(_03022_),
    .D(execution_unit_0.register_file_0.r8_15_ ),
    .Y(_02155_)
  );
  OAI21X1 _08779_ (
    .A(_02974_),
    .B(_03021_),
    .C(_02155_),
    .Y(_02156_)
  );
  AOI22X1 _08780_ (
    .A(execution_unit_0.register_file_0.r3_15_ ),
    .B(_03005_),
    .C(_03015_),
    .D(dbg_0.UNUSED_pc_15_ ),
    .Y(_02157_)
  );
  AOI22X1 _08781_ (
    .A(execution_unit_0.register_file_0.r10_15_ ),
    .B(_02992_),
    .C(_03011_),
    .D(execution_unit_0.register_file_0.r12_15_ ),
    .Y(_02158_)
  );
  NAND3X1 _08782_ (
    .A(_02154_),
    .B(_02157_),
    .C(_02158_),
    .Y(_02159_)
  );
  NOR2X1 _08783_ (
    .A(_02156_),
    .B(_02159_),
    .Y(_02160_)
  );
  AOI22X1 _08784_ (
    .A(execution_unit_0.register_file_0.r7_15_ ),
    .B(_02995_),
    .C(_03017_),
    .D(execution_unit_0.register_file_0.r9_15_ ),
    .Y(_02161_)
  );
  AOI22X1 _08785_ (
    .A(execution_unit_0.register_file_0.r13_15_ ),
    .B(_02990_),
    .C(_03007_),
    .D(execution_unit_0.register_file_0.r4_15_ ),
    .Y(_02162_)
  );
  NAND3X1 _08786_ (
    .A(_02153_),
    .B(_02161_),
    .C(_02162_),
    .Y(_02163_)
  );
  AOI21X1 _08787_ (
    .A(execution_unit_0.register_file_0.r14_15_ ),
    .B(_02997_),
    .C(_02163_),
    .Y(_02164_)
  );
  NAND2X1 _08788_ (
    .A(_02160_),
    .B(_02164_),
    .Y(execution_unit_0.reg_src_15_ )
  );
  XOR2X1 _08789_ (
    .A(_03302_),
    .B(execution_unit_0.reg_src_15_ ),
    .Y(_02165_)
  );
  OAI21X1 _08790_ (
    .A(execution_unit_0.register_file_0.r15_15_ ),
    .B(_03033_),
    .C(_03032_),
    .Y(_02166_)
  );
  INVX1 _08791_ (
    .A(_02166_),
    .Y(_02167_)
  );
  OAI21X1 _08792_ (
    .A(_03034_),
    .B(_02165_),
    .C(_02167_),
    .Y(_02168_)
  );
  OAI21X1 _08793_ (
    .A(_02989_),
    .B(_03032_),
    .C(_02168_),
    .Y(_02006_)
  );
  AND2X1 _08794_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_14_ ),
    .Y(_02169_)
  );
  NAND2X1 _08795_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_14_ ),
    .Y(_02170_)
  );
  AND2X1 _08796_ (
    .A(execution_unit_0.reg_incr ),
    .B(_02997_),
    .Y(_02171_)
  );
  NAND2X1 _08797_ (
    .A(execution_unit_0.reg_incr ),
    .B(_02997_),
    .Y(_02172_)
  );
  AOI21X1 _08798_ (
    .A(_03037_),
    .B(_02171_),
    .C(_02169_),
    .Y(_02173_)
  );
  OAI21X1 _08799_ (
    .A(execution_unit_0.register_file_0.r14_0_ ),
    .B(_02171_),
    .C(_02173_),
    .Y(_02174_)
  );
  OAI21X1 _08800_ (
    .A(_02955_),
    .B(_02170_),
    .C(_02174_),
    .Y(_01984_)
  );
  NOR2X1 _08801_ (
    .A(execution_unit_0.register_file_0.r14_1_ ),
    .B(_02171_),
    .Y(_02175_)
  );
  OAI21X1 _08802_ (
    .A(_03062_),
    .B(_02172_),
    .C(_02170_),
    .Y(_02176_)
  );
  OAI22X1 _08803_ (
    .A(_02956_),
    .B(_02170_),
    .C(_02175_),
    .D(_02176_),
    .Y(_01991_)
  );
  AOI21X1 _08804_ (
    .A(_03083_),
    .B(_02171_),
    .C(_02169_),
    .Y(_02177_)
  );
  OAI21X1 _08805_ (
    .A(execution_unit_0.register_file_0.r14_2_ ),
    .B(_02171_),
    .C(_02177_),
    .Y(_02178_)
  );
  OAI21X1 _08806_ (
    .A(_02959_),
    .B(_02170_),
    .C(_02178_),
    .Y(_01992_)
  );
  NOR2X1 _08807_ (
    .A(execution_unit_0.register_file_0.r14_3_ ),
    .B(_02171_),
    .Y(_02179_)
  );
  OAI21X1 _08808_ (
    .A(_03104_),
    .B(_02172_),
    .C(_02170_),
    .Y(_02180_)
  );
  OAI22X1 _08809_ (
    .A(_02962_),
    .B(_02170_),
    .C(_02179_),
    .D(_02180_),
    .Y(_01993_)
  );
  NOR2X1 _08810_ (
    .A(execution_unit_0.register_file_0.r14_4_ ),
    .B(_02171_),
    .Y(_02181_)
  );
  OAI21X1 _08811_ (
    .A(_03122_),
    .B(_02172_),
    .C(_02170_),
    .Y(_02182_)
  );
  OAI22X1 _08812_ (
    .A(_02965_),
    .B(_02170_),
    .C(_02181_),
    .D(_02182_),
    .Y(_01994_)
  );
  NOR2X1 _08813_ (
    .A(execution_unit_0.register_file_0.r14_5_ ),
    .B(_02171_),
    .Y(_02183_)
  );
  OAI21X1 _08814_ (
    .A(_03140_),
    .B(_02172_),
    .C(_02170_),
    .Y(_02184_)
  );
  OAI22X1 _08815_ (
    .A(_02966_),
    .B(_02170_),
    .C(_02183_),
    .D(_02184_),
    .Y(_01995_)
  );
  AOI21X1 _08816_ (
    .A(_03157_),
    .B(_02171_),
    .C(_02169_),
    .Y(_02185_)
  );
  OAI21X1 _08817_ (
    .A(execution_unit_0.register_file_0.r14_6_ ),
    .B(_02171_),
    .C(_02185_),
    .Y(_02186_)
  );
  OAI21X1 _08818_ (
    .A(_02967_),
    .B(_02170_),
    .C(_02186_),
    .Y(_01996_)
  );
  NOR2X1 _08819_ (
    .A(execution_unit_0.register_file_0.r14_7_ ),
    .B(_02171_),
    .Y(_02187_)
  );
  OAI21X1 _08820_ (
    .A(_03177_),
    .B(_02172_),
    .C(_02170_),
    .Y(_02188_)
  );
  OAI22X1 _08821_ (
    .A(_02968_),
    .B(_02170_),
    .C(_02187_),
    .D(_02188_),
    .Y(_01997_)
  );
  OAI21X1 _08822_ (
    .A(_03195_),
    .B(_02172_),
    .C(_02170_),
    .Y(_02189_)
  );
  INVX1 _08823_ (
    .A(_02189_),
    .Y(_02190_)
  );
  OAI21X1 _08824_ (
    .A(execution_unit_0.register_file_0.r14_8_ ),
    .B(_02171_),
    .C(_02190_),
    .Y(_02191_)
  );
  OAI21X1 _08825_ (
    .A(_02982_),
    .B(_02170_),
    .C(_02191_),
    .Y(_01998_)
  );
  OAI21X1 _08826_ (
    .A(_03212_),
    .B(_02172_),
    .C(_02170_),
    .Y(_02192_)
  );
  INVX1 _08827_ (
    .A(_02192_),
    .Y(_02193_)
  );
  OAI21X1 _08828_ (
    .A(execution_unit_0.register_file_0.r14_9_ ),
    .B(_02171_),
    .C(_02193_),
    .Y(_02194_)
  );
  OAI21X1 _08829_ (
    .A(_02983_),
    .B(_02170_),
    .C(_02194_),
    .Y(_01999_)
  );
  AOI21X1 _08830_ (
    .A(_03231_),
    .B(_02171_),
    .C(_02169_),
    .Y(_02195_)
  );
  OAI21X1 _08831_ (
    .A(execution_unit_0.register_file_0.r14_10_ ),
    .B(_02171_),
    .C(_02195_),
    .Y(_02196_)
  );
  OAI21X1 _08832_ (
    .A(_02984_),
    .B(_02170_),
    .C(_02196_),
    .Y(_01985_)
  );
  OAI21X1 _08833_ (
    .A(execution_unit_0.register_file_0.r14_11_ ),
    .B(_02171_),
    .C(_02170_),
    .Y(_02197_)
  );
  INVX1 _08834_ (
    .A(_02197_),
    .Y(_02198_)
  );
  OAI21X1 _08835_ (
    .A(_03249_),
    .B(_02172_),
    .C(_02198_),
    .Y(_02199_)
  );
  OAI21X1 _08836_ (
    .A(_02985_),
    .B(_02170_),
    .C(_02199_),
    .Y(_01986_)
  );
  OAI21X1 _08837_ (
    .A(execution_unit_0.register_file_0.r14_12_ ),
    .B(_02171_),
    .C(_02170_),
    .Y(_02200_)
  );
  INVX1 _08838_ (
    .A(_02200_),
    .Y(_02201_)
  );
  OAI21X1 _08839_ (
    .A(_03267_),
    .B(_02172_),
    .C(_02201_),
    .Y(_02202_)
  );
  OAI21X1 _08840_ (
    .A(_02986_),
    .B(_02170_),
    .C(_02202_),
    .Y(_01987_)
  );
  OAI21X1 _08841_ (
    .A(execution_unit_0.register_file_0.r14_13_ ),
    .B(_02171_),
    .C(_02170_),
    .Y(_02203_)
  );
  INVX1 _08842_ (
    .A(_02203_),
    .Y(_02204_)
  );
  OAI21X1 _08843_ (
    .A(_03285_),
    .B(_02172_),
    .C(_02204_),
    .Y(_02205_)
  );
  OAI21X1 _08844_ (
    .A(_02987_),
    .B(_02170_),
    .C(_02205_),
    .Y(_01988_)
  );
  OAI21X1 _08845_ (
    .A(execution_unit_0.register_file_0.r14_14_ ),
    .B(_02171_),
    .C(_02170_),
    .Y(_02206_)
  );
  INVX1 _08846_ (
    .A(_02206_),
    .Y(_02207_)
  );
  OAI21X1 _08847_ (
    .A(_03303_),
    .B(_02172_),
    .C(_02207_),
    .Y(_02208_)
  );
  OAI21X1 _08848_ (
    .A(_02988_),
    .B(_02170_),
    .C(_02208_),
    .Y(_01989_)
  );
  OAI21X1 _08849_ (
    .A(execution_unit_0.register_file_0.r14_15_ ),
    .B(_02171_),
    .C(_02170_),
    .Y(_02209_)
  );
  INVX1 _08850_ (
    .A(_02209_),
    .Y(_02210_)
  );
  OAI21X1 _08851_ (
    .A(_02165_),
    .B(_02172_),
    .C(_02210_),
    .Y(_02211_)
  );
  OAI21X1 _08852_ (
    .A(_02989_),
    .B(_02170_),
    .C(_02211_),
    .Y(_01990_)
  );
  AND2X1 _08853_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_13_ ),
    .Y(_02212_)
  );
  NAND2X1 _08854_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_13_ ),
    .Y(_02213_)
  );
  AND2X1 _08855_ (
    .A(execution_unit_0.reg_incr ),
    .B(_02990_),
    .Y(_02214_)
  );
  NAND2X1 _08856_ (
    .A(execution_unit_0.reg_incr ),
    .B(_02990_),
    .Y(_02215_)
  );
  AOI21X1 _08857_ (
    .A(_03037_),
    .B(_02214_),
    .C(_02212_),
    .Y(_02216_)
  );
  OAI21X1 _08858_ (
    .A(execution_unit_0.register_file_0.r13_0_ ),
    .B(_02214_),
    .C(_02216_),
    .Y(_02217_)
  );
  OAI21X1 _08859_ (
    .A(_02955_),
    .B(_02213_),
    .C(_02217_),
    .Y(_01968_)
  );
  NOR2X1 _08860_ (
    .A(execution_unit_0.register_file_0.r13_1_ ),
    .B(_02214_),
    .Y(_02218_)
  );
  OAI21X1 _08861_ (
    .A(_03062_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02219_)
  );
  OAI22X1 _08862_ (
    .A(_02956_),
    .B(_02213_),
    .C(_02218_),
    .D(_02219_),
    .Y(_01975_)
  );
  AND2X1 _08863_ (
    .A(_03083_),
    .B(_02214_),
    .Y(_02220_)
  );
  OAI21X1 _08864_ (
    .A(execution_unit_0.register_file_0.r13_2_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02221_)
  );
  OAI22X1 _08865_ (
    .A(_02959_),
    .B(_02213_),
    .C(_02220_),
    .D(_02221_),
    .Y(_01976_)
  );
  NOR2X1 _08866_ (
    .A(execution_unit_0.register_file_0.r13_3_ ),
    .B(_02214_),
    .Y(_02222_)
  );
  OAI21X1 _08867_ (
    .A(_03104_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02223_)
  );
  OAI22X1 _08868_ (
    .A(_02962_),
    .B(_02213_),
    .C(_02222_),
    .D(_02223_),
    .Y(_01977_)
  );
  NOR2X1 _08869_ (
    .A(execution_unit_0.register_file_0.r13_4_ ),
    .B(_02214_),
    .Y(_02224_)
  );
  OAI21X1 _08870_ (
    .A(_03122_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02225_)
  );
  OAI22X1 _08871_ (
    .A(_02965_),
    .B(_02213_),
    .C(_02224_),
    .D(_02225_),
    .Y(_01978_)
  );
  NOR2X1 _08872_ (
    .A(execution_unit_0.register_file_0.r13_5_ ),
    .B(_02214_),
    .Y(_02226_)
  );
  OAI21X1 _08873_ (
    .A(_03140_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02227_)
  );
  OAI22X1 _08874_ (
    .A(_02966_),
    .B(_02213_),
    .C(_02226_),
    .D(_02227_),
    .Y(_01979_)
  );
  AOI21X1 _08875_ (
    .A(_03157_),
    .B(_02214_),
    .C(_02212_),
    .Y(_02228_)
  );
  OAI21X1 _08876_ (
    .A(execution_unit_0.register_file_0.r13_6_ ),
    .B(_02214_),
    .C(_02228_),
    .Y(_02229_)
  );
  OAI21X1 _08877_ (
    .A(_02967_),
    .B(_02213_),
    .C(_02229_),
    .Y(_01980_)
  );
  NOR2X1 _08878_ (
    .A(execution_unit_0.register_file_0.r13_7_ ),
    .B(_02214_),
    .Y(_02230_)
  );
  OAI21X1 _08879_ (
    .A(_03177_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02231_)
  );
  OAI22X1 _08880_ (
    .A(_02968_),
    .B(_02213_),
    .C(_02230_),
    .D(_02231_),
    .Y(_01981_)
  );
  OAI21X1 _08881_ (
    .A(_03195_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02232_)
  );
  INVX1 _08882_ (
    .A(_02232_),
    .Y(_02233_)
  );
  OAI21X1 _08883_ (
    .A(execution_unit_0.register_file_0.r13_8_ ),
    .B(_02214_),
    .C(_02233_),
    .Y(_02234_)
  );
  OAI21X1 _08884_ (
    .A(_02982_),
    .B(_02213_),
    .C(_02234_),
    .Y(_01982_)
  );
  OAI21X1 _08885_ (
    .A(_03212_),
    .B(_02215_),
    .C(_02213_),
    .Y(_02235_)
  );
  INVX1 _08886_ (
    .A(_02235_),
    .Y(_02236_)
  );
  OAI21X1 _08887_ (
    .A(execution_unit_0.register_file_0.r13_9_ ),
    .B(_02214_),
    .C(_02236_),
    .Y(_02237_)
  );
  OAI21X1 _08888_ (
    .A(_02983_),
    .B(_02213_),
    .C(_02237_),
    .Y(_01983_)
  );
  AOI21X1 _08889_ (
    .A(_03231_),
    .B(_02214_),
    .C(_02212_),
    .Y(_02238_)
  );
  OAI21X1 _08890_ (
    .A(execution_unit_0.register_file_0.r13_10_ ),
    .B(_02214_),
    .C(_02238_),
    .Y(_02239_)
  );
  OAI21X1 _08891_ (
    .A(_02984_),
    .B(_02213_),
    .C(_02239_),
    .Y(_01969_)
  );
  OAI21X1 _08892_ (
    .A(execution_unit_0.register_file_0.r13_11_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02240_)
  );
  INVX1 _08893_ (
    .A(_02240_),
    .Y(_02241_)
  );
  OAI21X1 _08894_ (
    .A(_03249_),
    .B(_02215_),
    .C(_02241_),
    .Y(_02242_)
  );
  OAI21X1 _08895_ (
    .A(_02985_),
    .B(_02213_),
    .C(_02242_),
    .Y(_01970_)
  );
  OAI21X1 _08896_ (
    .A(execution_unit_0.register_file_0.r13_12_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02243_)
  );
  INVX1 _08897_ (
    .A(_02243_),
    .Y(_02244_)
  );
  OAI21X1 _08898_ (
    .A(_03267_),
    .B(_02215_),
    .C(_02244_),
    .Y(_02245_)
  );
  OAI21X1 _08899_ (
    .A(_02986_),
    .B(_02213_),
    .C(_02245_),
    .Y(_01971_)
  );
  OAI21X1 _08900_ (
    .A(execution_unit_0.register_file_0.r13_13_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02246_)
  );
  INVX1 _08901_ (
    .A(_02246_),
    .Y(_02247_)
  );
  OAI21X1 _08902_ (
    .A(_03285_),
    .B(_02215_),
    .C(_02247_),
    .Y(_02248_)
  );
  OAI21X1 _08903_ (
    .A(_02987_),
    .B(_02213_),
    .C(_02248_),
    .Y(_01972_)
  );
  OAI21X1 _08904_ (
    .A(execution_unit_0.register_file_0.r13_14_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02249_)
  );
  INVX1 _08905_ (
    .A(_02249_),
    .Y(_02250_)
  );
  OAI21X1 _08906_ (
    .A(_03303_),
    .B(_02215_),
    .C(_02250_),
    .Y(_02251_)
  );
  OAI21X1 _08907_ (
    .A(_02988_),
    .B(_02213_),
    .C(_02251_),
    .Y(_01973_)
  );
  OAI21X1 _08908_ (
    .A(execution_unit_0.register_file_0.r13_15_ ),
    .B(_02214_),
    .C(_02213_),
    .Y(_02252_)
  );
  INVX1 _08909_ (
    .A(_02252_),
    .Y(_02253_)
  );
  OAI21X1 _08910_ (
    .A(_02165_),
    .B(_02215_),
    .C(_02253_),
    .Y(_02254_)
  );
  OAI21X1 _08911_ (
    .A(_02989_),
    .B(_02213_),
    .C(_02254_),
    .Y(_01974_)
  );
  AND2X1 _08912_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_12_ ),
    .Y(_02255_)
  );
  NAND2X1 _08913_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_12_ ),
    .Y(_02256_)
  );
  AND2X1 _08914_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03011_),
    .Y(_02257_)
  );
  NAND2X1 _08915_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03011_),
    .Y(_02258_)
  );
  AOI21X1 _08916_ (
    .A(_03037_),
    .B(_02257_),
    .C(_02255_),
    .Y(_02259_)
  );
  OAI21X1 _08917_ (
    .A(execution_unit_0.register_file_0.r12_0_ ),
    .B(_02257_),
    .C(_02259_),
    .Y(_02260_)
  );
  OAI21X1 _08918_ (
    .A(_02955_),
    .B(_02256_),
    .C(_02260_),
    .Y(_01952_)
  );
  NOR2X1 _08919_ (
    .A(execution_unit_0.register_file_0.r12_1_ ),
    .B(_02257_),
    .Y(_02261_)
  );
  OAI21X1 _08920_ (
    .A(_03062_),
    .B(_02258_),
    .C(_02256_),
    .Y(_02262_)
  );
  OAI22X1 _08921_ (
    .A(_02956_),
    .B(_02256_),
    .C(_02261_),
    .D(_02262_),
    .Y(_01959_)
  );
  AOI21X1 _08922_ (
    .A(_03083_),
    .B(_02257_),
    .C(_02255_),
    .Y(_02263_)
  );
  OAI21X1 _08923_ (
    .A(execution_unit_0.register_file_0.r12_2_ ),
    .B(_02257_),
    .C(_02263_),
    .Y(_02264_)
  );
  OAI21X1 _08924_ (
    .A(_02959_),
    .B(_02256_),
    .C(_02264_),
    .Y(_01960_)
  );
  NOR2X1 _08925_ (
    .A(execution_unit_0.register_file_0.r12_3_ ),
    .B(_02257_),
    .Y(_02265_)
  );
  OAI21X1 _08926_ (
    .A(_03104_),
    .B(_02258_),
    .C(_02256_),
    .Y(_02266_)
  );
  OAI22X1 _08927_ (
    .A(_02962_),
    .B(_02256_),
    .C(_02265_),
    .D(_02266_),
    .Y(_01961_)
  );
  NOR2X1 _08928_ (
    .A(execution_unit_0.register_file_0.r12_4_ ),
    .B(_02257_),
    .Y(_02267_)
  );
  OAI21X1 _08929_ (
    .A(_03122_),
    .B(_02258_),
    .C(_02256_),
    .Y(_02268_)
  );
  OAI22X1 _08930_ (
    .A(_02965_),
    .B(_02256_),
    .C(_02267_),
    .D(_02268_),
    .Y(_01962_)
  );
  NOR2X1 _08931_ (
    .A(execution_unit_0.register_file_0.r12_5_ ),
    .B(_02257_),
    .Y(_02269_)
  );
  OAI21X1 _08932_ (
    .A(_03140_),
    .B(_02258_),
    .C(_02256_),
    .Y(_02270_)
  );
  OAI22X1 _08933_ (
    .A(_02966_),
    .B(_02256_),
    .C(_02269_),
    .D(_02270_),
    .Y(_01963_)
  );
  AOI21X1 _08934_ (
    .A(_03157_),
    .B(_02257_),
    .C(_02255_),
    .Y(_02271_)
  );
  OAI21X1 _08935_ (
    .A(execution_unit_0.register_file_0.r12_6_ ),
    .B(_02257_),
    .C(_02271_),
    .Y(_02272_)
  );
  OAI21X1 _08936_ (
    .A(_02967_),
    .B(_02256_),
    .C(_02272_),
    .Y(_01964_)
  );
  NOR2X1 _08937_ (
    .A(execution_unit_0.register_file_0.r12_7_ ),
    .B(_02257_),
    .Y(_02273_)
  );
  OAI21X1 _08938_ (
    .A(_03177_),
    .B(_02258_),
    .C(_02256_),
    .Y(_02274_)
  );
  OAI22X1 _08939_ (
    .A(_02968_),
    .B(_02256_),
    .C(_02273_),
    .D(_02274_),
    .Y(_01965_)
  );
  OAI21X1 _08940_ (
    .A(_03195_),
    .B(_02258_),
    .C(_02256_),
    .Y(_02275_)
  );
  INVX1 _08941_ (
    .A(_02275_),
    .Y(_02276_)
  );
  OAI21X1 _08942_ (
    .A(execution_unit_0.register_file_0.r12_8_ ),
    .B(_02257_),
    .C(_02276_),
    .Y(_02277_)
  );
  OAI21X1 _08943_ (
    .A(_02982_),
    .B(_02256_),
    .C(_02277_),
    .Y(_01966_)
  );
  OAI21X1 _08944_ (
    .A(_03212_),
    .B(_02258_),
    .C(_02256_),
    .Y(_02278_)
  );
  INVX1 _08945_ (
    .A(_02278_),
    .Y(_02279_)
  );
  OAI21X1 _08946_ (
    .A(execution_unit_0.register_file_0.r12_9_ ),
    .B(_02257_),
    .C(_02279_),
    .Y(_02280_)
  );
  OAI21X1 _08947_ (
    .A(_02983_),
    .B(_02256_),
    .C(_02280_),
    .Y(_01967_)
  );
  AOI21X1 _08948_ (
    .A(_03231_),
    .B(_02257_),
    .C(_02255_),
    .Y(_02281_)
  );
  OAI21X1 _08949_ (
    .A(execution_unit_0.register_file_0.r12_10_ ),
    .B(_02257_),
    .C(_02281_),
    .Y(_02282_)
  );
  OAI21X1 _08950_ (
    .A(_02984_),
    .B(_02256_),
    .C(_02282_),
    .Y(_01953_)
  );
  OAI21X1 _08951_ (
    .A(execution_unit_0.register_file_0.r12_11_ ),
    .B(_02257_),
    .C(_02256_),
    .Y(_02283_)
  );
  INVX1 _08952_ (
    .A(_02283_),
    .Y(_02284_)
  );
  OAI21X1 _08953_ (
    .A(_03249_),
    .B(_02258_),
    .C(_02284_),
    .Y(_02285_)
  );
  OAI21X1 _08954_ (
    .A(_02985_),
    .B(_02256_),
    .C(_02285_),
    .Y(_01954_)
  );
  OAI21X1 _08955_ (
    .A(execution_unit_0.register_file_0.r12_12_ ),
    .B(_02257_),
    .C(_02256_),
    .Y(_02286_)
  );
  INVX1 _08956_ (
    .A(_02286_),
    .Y(_02287_)
  );
  OAI21X1 _08957_ (
    .A(_03267_),
    .B(_02258_),
    .C(_02287_),
    .Y(_02288_)
  );
  OAI21X1 _08958_ (
    .A(_02986_),
    .B(_02256_),
    .C(_02288_),
    .Y(_01955_)
  );
  OAI21X1 _08959_ (
    .A(execution_unit_0.register_file_0.r12_13_ ),
    .B(_02257_),
    .C(_02256_),
    .Y(_02289_)
  );
  INVX1 _08960_ (
    .A(_02289_),
    .Y(_02290_)
  );
  OAI21X1 _08961_ (
    .A(_03285_),
    .B(_02258_),
    .C(_02290_),
    .Y(_02291_)
  );
  OAI21X1 _08962_ (
    .A(_02987_),
    .B(_02256_),
    .C(_02291_),
    .Y(_01956_)
  );
  OAI21X1 _08963_ (
    .A(execution_unit_0.register_file_0.r12_14_ ),
    .B(_02257_),
    .C(_02256_),
    .Y(_02292_)
  );
  INVX1 _08964_ (
    .A(_02292_),
    .Y(_02293_)
  );
  OAI21X1 _08965_ (
    .A(_03303_),
    .B(_02258_),
    .C(_02293_),
    .Y(_02294_)
  );
  OAI21X1 _08966_ (
    .A(_02988_),
    .B(_02256_),
    .C(_02294_),
    .Y(_01957_)
  );
  OAI21X1 _08967_ (
    .A(execution_unit_0.register_file_0.r12_15_ ),
    .B(_02257_),
    .C(_02256_),
    .Y(_02295_)
  );
  INVX1 _08968_ (
    .A(_02295_),
    .Y(_02296_)
  );
  OAI21X1 _08969_ (
    .A(_02165_),
    .B(_02258_),
    .C(_02296_),
    .Y(_02297_)
  );
  OAI21X1 _08970_ (
    .A(_02989_),
    .B(_02256_),
    .C(_02297_),
    .Y(_01958_)
  );
  AND2X1 _08971_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_11_ ),
    .Y(_02298_)
  );
  NAND2X1 _08972_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_11_ ),
    .Y(_02299_)
  );
  AND2X1 _08973_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03009_),
    .Y(_02300_)
  );
  NAND2X1 _08974_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03009_),
    .Y(_02301_)
  );
  AOI21X1 _08975_ (
    .A(_03037_),
    .B(_02300_),
    .C(_02298_),
    .Y(_02302_)
  );
  OAI21X1 _08976_ (
    .A(execution_unit_0.register_file_0.r11_0_ ),
    .B(_02300_),
    .C(_02302_),
    .Y(_02303_)
  );
  OAI21X1 _08977_ (
    .A(_02955_),
    .B(_02299_),
    .C(_02303_),
    .Y(_01936_)
  );
  NOR2X1 _08978_ (
    .A(execution_unit_0.register_file_0.r11_1_ ),
    .B(_02300_),
    .Y(_02304_)
  );
  OAI21X1 _08979_ (
    .A(_03062_),
    .B(_02301_),
    .C(_02299_),
    .Y(_02305_)
  );
  OAI22X1 _08980_ (
    .A(_02956_),
    .B(_02299_),
    .C(_02304_),
    .D(_02305_),
    .Y(_01943_)
  );
  AOI21X1 _08981_ (
    .A(_03083_),
    .B(_02300_),
    .C(_02298_),
    .Y(_02306_)
  );
  OAI21X1 _08982_ (
    .A(execution_unit_0.register_file_0.r11_2_ ),
    .B(_02300_),
    .C(_02306_),
    .Y(_02307_)
  );
  OAI21X1 _08983_ (
    .A(_02959_),
    .B(_02299_),
    .C(_02307_),
    .Y(_01944_)
  );
  NOR2X1 _08984_ (
    .A(execution_unit_0.register_file_0.r11_3_ ),
    .B(_02300_),
    .Y(_02308_)
  );
  OAI21X1 _08985_ (
    .A(_03104_),
    .B(_02301_),
    .C(_02299_),
    .Y(_02309_)
  );
  OAI22X1 _08986_ (
    .A(_02962_),
    .B(_02299_),
    .C(_02308_),
    .D(_02309_),
    .Y(_01945_)
  );
  NOR2X1 _08987_ (
    .A(execution_unit_0.register_file_0.r11_4_ ),
    .B(_02300_),
    .Y(_02310_)
  );
  OAI21X1 _08988_ (
    .A(_03122_),
    .B(_02301_),
    .C(_02299_),
    .Y(_02311_)
  );
  OAI22X1 _08989_ (
    .A(_02965_),
    .B(_02299_),
    .C(_02310_),
    .D(_02311_),
    .Y(_01946_)
  );
  NOR2X1 _08990_ (
    .A(execution_unit_0.register_file_0.r11_5_ ),
    .B(_02300_),
    .Y(_02312_)
  );
  OAI21X1 _08991_ (
    .A(_03140_),
    .B(_02301_),
    .C(_02299_),
    .Y(_02313_)
  );
  OAI22X1 _08992_ (
    .A(_02966_),
    .B(_02299_),
    .C(_02312_),
    .D(_02313_),
    .Y(_01947_)
  );
  AOI21X1 _08993_ (
    .A(_03157_),
    .B(_02300_),
    .C(_02298_),
    .Y(_02314_)
  );
  OAI21X1 _08994_ (
    .A(execution_unit_0.register_file_0.r11_6_ ),
    .B(_02300_),
    .C(_02314_),
    .Y(_02315_)
  );
  OAI21X1 _08995_ (
    .A(_02967_),
    .B(_02299_),
    .C(_02315_),
    .Y(_01948_)
  );
  NOR2X1 _08996_ (
    .A(execution_unit_0.register_file_0.r11_7_ ),
    .B(_02300_),
    .Y(_02316_)
  );
  OAI21X1 _08997_ (
    .A(_03177_),
    .B(_02301_),
    .C(_02299_),
    .Y(_02317_)
  );
  OAI22X1 _08998_ (
    .A(_02968_),
    .B(_02299_),
    .C(_02316_),
    .D(_02317_),
    .Y(_01949_)
  );
  OAI21X1 _08999_ (
    .A(_03195_),
    .B(_02301_),
    .C(_02299_),
    .Y(_02318_)
  );
  INVX1 _09000_ (
    .A(_02318_),
    .Y(_02319_)
  );
  OAI21X1 _09001_ (
    .A(execution_unit_0.register_file_0.r11_8_ ),
    .B(_02300_),
    .C(_02319_),
    .Y(_02320_)
  );
  OAI21X1 _09002_ (
    .A(_02982_),
    .B(_02299_),
    .C(_02320_),
    .Y(_01950_)
  );
  OAI21X1 _09003_ (
    .A(_03212_),
    .B(_02301_),
    .C(_02299_),
    .Y(_02321_)
  );
  INVX1 _09004_ (
    .A(_02321_),
    .Y(_02322_)
  );
  OAI21X1 _09005_ (
    .A(execution_unit_0.register_file_0.r11_9_ ),
    .B(_02300_),
    .C(_02322_),
    .Y(_02323_)
  );
  OAI21X1 _09006_ (
    .A(_02983_),
    .B(_02299_),
    .C(_02323_),
    .Y(_01951_)
  );
  AOI21X1 _09007_ (
    .A(_03231_),
    .B(_02300_),
    .C(_02298_),
    .Y(_02324_)
  );
  OAI21X1 _09008_ (
    .A(execution_unit_0.register_file_0.r11_10_ ),
    .B(_02300_),
    .C(_02324_),
    .Y(_02325_)
  );
  OAI21X1 _09009_ (
    .A(_02984_),
    .B(_02299_),
    .C(_02325_),
    .Y(_01937_)
  );
  OAI21X1 _09010_ (
    .A(execution_unit_0.register_file_0.r11_11_ ),
    .B(_02300_),
    .C(_02299_),
    .Y(_02326_)
  );
  INVX1 _09011_ (
    .A(_02326_),
    .Y(_02327_)
  );
  OAI21X1 _09012_ (
    .A(_03249_),
    .B(_02301_),
    .C(_02327_),
    .Y(_02328_)
  );
  OAI21X1 _09013_ (
    .A(_02985_),
    .B(_02299_),
    .C(_02328_),
    .Y(_01938_)
  );
  OAI21X1 _09014_ (
    .A(execution_unit_0.register_file_0.r11_12_ ),
    .B(_02300_),
    .C(_02299_),
    .Y(_02329_)
  );
  INVX1 _09015_ (
    .A(_02329_),
    .Y(_02330_)
  );
  OAI21X1 _09016_ (
    .A(_03267_),
    .B(_02301_),
    .C(_02330_),
    .Y(_02331_)
  );
  OAI21X1 _09017_ (
    .A(_02986_),
    .B(_02299_),
    .C(_02331_),
    .Y(_01939_)
  );
  OAI21X1 _09018_ (
    .A(execution_unit_0.register_file_0.r11_13_ ),
    .B(_02300_),
    .C(_02299_),
    .Y(_02332_)
  );
  INVX1 _09019_ (
    .A(_02332_),
    .Y(_02333_)
  );
  OAI21X1 _09020_ (
    .A(_03285_),
    .B(_02301_),
    .C(_02333_),
    .Y(_02334_)
  );
  OAI21X1 _09021_ (
    .A(_02987_),
    .B(_02299_),
    .C(_02334_),
    .Y(_01940_)
  );
  OAI21X1 _09022_ (
    .A(execution_unit_0.register_file_0.r11_14_ ),
    .B(_02300_),
    .C(_02299_),
    .Y(_02335_)
  );
  INVX1 _09023_ (
    .A(_02335_),
    .Y(_02336_)
  );
  OAI21X1 _09024_ (
    .A(_03303_),
    .B(_02301_),
    .C(_02336_),
    .Y(_02337_)
  );
  OAI21X1 _09025_ (
    .A(_02988_),
    .B(_02299_),
    .C(_02337_),
    .Y(_01941_)
  );
  OAI21X1 _09026_ (
    .A(execution_unit_0.register_file_0.r11_15_ ),
    .B(_02300_),
    .C(_02299_),
    .Y(_02338_)
  );
  INVX1 _09027_ (
    .A(_02338_),
    .Y(_02339_)
  );
  OAI21X1 _09028_ (
    .A(_02165_),
    .B(_02301_),
    .C(_02339_),
    .Y(_02340_)
  );
  OAI21X1 _09029_ (
    .A(_02989_),
    .B(_02299_),
    .C(_02340_),
    .Y(_01942_)
  );
  AND2X1 _09030_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_10_ ),
    .Y(_02341_)
  );
  NAND2X1 _09031_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_10_ ),
    .Y(_02342_)
  );
  AND2X1 _09032_ (
    .A(execution_unit_0.reg_incr ),
    .B(_02992_),
    .Y(_02343_)
  );
  NAND2X1 _09033_ (
    .A(execution_unit_0.reg_incr ),
    .B(_02992_),
    .Y(_02344_)
  );
  AOI21X1 _09034_ (
    .A(_03037_),
    .B(_02343_),
    .C(_02341_),
    .Y(_02345_)
  );
  OAI21X1 _09035_ (
    .A(execution_unit_0.register_file_0.r10_0_ ),
    .B(_02343_),
    .C(_02345_),
    .Y(_02346_)
  );
  OAI21X1 _09036_ (
    .A(_02955_),
    .B(_02342_),
    .C(_02346_),
    .Y(_01920_)
  );
  NOR2X1 _09037_ (
    .A(execution_unit_0.register_file_0.r10_1_ ),
    .B(_02343_),
    .Y(_02347_)
  );
  OAI21X1 _09038_ (
    .A(_03062_),
    .B(_02344_),
    .C(_02342_),
    .Y(_02348_)
  );
  OAI22X1 _09039_ (
    .A(_02956_),
    .B(_02342_),
    .C(_02347_),
    .D(_02348_),
    .Y(_01927_)
  );
  AOI21X1 _09040_ (
    .A(_03083_),
    .B(_02343_),
    .C(_02341_),
    .Y(_02349_)
  );
  OAI21X1 _09041_ (
    .A(execution_unit_0.register_file_0.r10_2_ ),
    .B(_02343_),
    .C(_02349_),
    .Y(_02350_)
  );
  OAI21X1 _09042_ (
    .A(_02959_),
    .B(_02342_),
    .C(_02350_),
    .Y(_01928_)
  );
  NOR2X1 _09043_ (
    .A(execution_unit_0.register_file_0.r10_3_ ),
    .B(_02343_),
    .Y(_02351_)
  );
  OAI21X1 _09044_ (
    .A(_03104_),
    .B(_02344_),
    .C(_02342_),
    .Y(_02352_)
  );
  OAI22X1 _09045_ (
    .A(_02962_),
    .B(_02342_),
    .C(_02351_),
    .D(_02352_),
    .Y(_01929_)
  );
  NOR2X1 _09046_ (
    .A(execution_unit_0.register_file_0.r10_4_ ),
    .B(_02343_),
    .Y(_02353_)
  );
  OAI21X1 _09047_ (
    .A(_03122_),
    .B(_02344_),
    .C(_02342_),
    .Y(_02354_)
  );
  OAI22X1 _09048_ (
    .A(_02965_),
    .B(_02342_),
    .C(_02353_),
    .D(_02354_),
    .Y(_01930_)
  );
  NOR2X1 _09049_ (
    .A(execution_unit_0.register_file_0.r10_5_ ),
    .B(_02343_),
    .Y(_02355_)
  );
  OAI21X1 _09050_ (
    .A(_03140_),
    .B(_02344_),
    .C(_02342_),
    .Y(_02356_)
  );
  OAI22X1 _09051_ (
    .A(_02966_),
    .B(_02342_),
    .C(_02355_),
    .D(_02356_),
    .Y(_01931_)
  );
  AOI21X1 _09052_ (
    .A(_03157_),
    .B(_02343_),
    .C(_02341_),
    .Y(_02357_)
  );
  OAI21X1 _09053_ (
    .A(execution_unit_0.register_file_0.r10_6_ ),
    .B(_02343_),
    .C(_02357_),
    .Y(_02358_)
  );
  OAI21X1 _09054_ (
    .A(_02967_),
    .B(_02342_),
    .C(_02358_),
    .Y(_01932_)
  );
  NOR2X1 _09055_ (
    .A(execution_unit_0.register_file_0.r10_7_ ),
    .B(_02343_),
    .Y(_02359_)
  );
  OAI21X1 _09056_ (
    .A(_03177_),
    .B(_02344_),
    .C(_02342_),
    .Y(_02360_)
  );
  OAI22X1 _09057_ (
    .A(_02968_),
    .B(_02342_),
    .C(_02359_),
    .D(_02360_),
    .Y(_01933_)
  );
  OAI21X1 _09058_ (
    .A(_03195_),
    .B(_02344_),
    .C(_02342_),
    .Y(_02361_)
  );
  INVX1 _09059_ (
    .A(_02361_),
    .Y(_02362_)
  );
  OAI21X1 _09060_ (
    .A(execution_unit_0.register_file_0.r10_8_ ),
    .B(_02343_),
    .C(_02362_),
    .Y(_02363_)
  );
  OAI21X1 _09061_ (
    .A(_02982_),
    .B(_02342_),
    .C(_02363_),
    .Y(_01934_)
  );
  OAI21X1 _09062_ (
    .A(_03212_),
    .B(_02344_),
    .C(_02342_),
    .Y(_02364_)
  );
  INVX1 _09063_ (
    .A(_02364_),
    .Y(_02365_)
  );
  OAI21X1 _09064_ (
    .A(execution_unit_0.register_file_0.r10_9_ ),
    .B(_02343_),
    .C(_02365_),
    .Y(_02366_)
  );
  OAI21X1 _09065_ (
    .A(_02983_),
    .B(_02342_),
    .C(_02366_),
    .Y(_01935_)
  );
  AOI21X1 _09066_ (
    .A(_03231_),
    .B(_02343_),
    .C(_02341_),
    .Y(_02367_)
  );
  OAI21X1 _09067_ (
    .A(execution_unit_0.register_file_0.r10_10_ ),
    .B(_02343_),
    .C(_02367_),
    .Y(_02368_)
  );
  OAI21X1 _09068_ (
    .A(_02984_),
    .B(_02342_),
    .C(_02368_),
    .Y(_01921_)
  );
  OAI21X1 _09069_ (
    .A(execution_unit_0.register_file_0.r10_11_ ),
    .B(_02343_),
    .C(_02342_),
    .Y(_02369_)
  );
  INVX1 _09070_ (
    .A(_02369_),
    .Y(_02370_)
  );
  OAI21X1 _09071_ (
    .A(_03249_),
    .B(_02344_),
    .C(_02370_),
    .Y(_02371_)
  );
  OAI21X1 _09072_ (
    .A(_02985_),
    .B(_02342_),
    .C(_02371_),
    .Y(_01922_)
  );
  OAI21X1 _09073_ (
    .A(execution_unit_0.register_file_0.r10_12_ ),
    .B(_02343_),
    .C(_02342_),
    .Y(_02372_)
  );
  INVX1 _09074_ (
    .A(_02372_),
    .Y(_02373_)
  );
  OAI21X1 _09075_ (
    .A(_03267_),
    .B(_02344_),
    .C(_02373_),
    .Y(_02374_)
  );
  OAI21X1 _09076_ (
    .A(_02986_),
    .B(_02342_),
    .C(_02374_),
    .Y(_01923_)
  );
  OAI21X1 _09077_ (
    .A(execution_unit_0.register_file_0.r10_13_ ),
    .B(_02343_),
    .C(_02342_),
    .Y(_02375_)
  );
  INVX1 _09078_ (
    .A(_02375_),
    .Y(_02376_)
  );
  OAI21X1 _09079_ (
    .A(_03285_),
    .B(_02344_),
    .C(_02376_),
    .Y(_02377_)
  );
  OAI21X1 _09080_ (
    .A(_02987_),
    .B(_02342_),
    .C(_02377_),
    .Y(_01924_)
  );
  OAI21X1 _09081_ (
    .A(execution_unit_0.register_file_0.r10_14_ ),
    .B(_02343_),
    .C(_02342_),
    .Y(_02378_)
  );
  INVX1 _09082_ (
    .A(_02378_),
    .Y(_02379_)
  );
  OAI21X1 _09083_ (
    .A(_03303_),
    .B(_02344_),
    .C(_02379_),
    .Y(_02380_)
  );
  OAI21X1 _09084_ (
    .A(_02988_),
    .B(_02342_),
    .C(_02380_),
    .Y(_01925_)
  );
  OAI21X1 _09085_ (
    .A(execution_unit_0.register_file_0.r10_15_ ),
    .B(_02343_),
    .C(_02342_),
    .Y(_02381_)
  );
  INVX1 _09086_ (
    .A(_02381_),
    .Y(_02382_)
  );
  OAI21X1 _09087_ (
    .A(_02165_),
    .B(_02344_),
    .C(_02382_),
    .Y(_02383_)
  );
  OAI21X1 _09088_ (
    .A(_02989_),
    .B(_02342_),
    .C(_02383_),
    .Y(_01926_)
  );
  AND2X1 _09089_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_9_ ),
    .Y(_02384_)
  );
  NAND2X1 _09090_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_9_ ),
    .Y(_02385_)
  );
  AND2X1 _09091_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03017_),
    .Y(_02386_)
  );
  NAND2X1 _09092_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03017_),
    .Y(_02387_)
  );
  AOI21X1 _09093_ (
    .A(_03037_),
    .B(_02386_),
    .C(_02384_),
    .Y(_02388_)
  );
  OAI21X1 _09094_ (
    .A(execution_unit_0.register_file_0.r9_0_ ),
    .B(_02386_),
    .C(_02388_),
    .Y(_02389_)
  );
  OAI21X1 _09095_ (
    .A(_02955_),
    .B(_02385_),
    .C(_02389_),
    .Y(_02136_)
  );
  NOR2X1 _09096_ (
    .A(execution_unit_0.register_file_0.r9_1_ ),
    .B(_02386_),
    .Y(_02390_)
  );
  OAI21X1 _09097_ (
    .A(_03062_),
    .B(_02387_),
    .C(_02385_),
    .Y(_02391_)
  );
  OAI22X1 _09098_ (
    .A(_02956_),
    .B(_02385_),
    .C(_02390_),
    .D(_02391_),
    .Y(_02143_)
  );
  AOI21X1 _09099_ (
    .A(_03083_),
    .B(_02386_),
    .C(_02384_),
    .Y(_02392_)
  );
  OAI21X1 _09100_ (
    .A(execution_unit_0.register_file_0.r9_2_ ),
    .B(_02386_),
    .C(_02392_),
    .Y(_02393_)
  );
  OAI21X1 _09101_ (
    .A(_02959_),
    .B(_02385_),
    .C(_02393_),
    .Y(_02144_)
  );
  NOR2X1 _09102_ (
    .A(execution_unit_0.register_file_0.r9_3_ ),
    .B(_02386_),
    .Y(_02394_)
  );
  OAI21X1 _09103_ (
    .A(_03104_),
    .B(_02387_),
    .C(_02385_),
    .Y(_02395_)
  );
  OAI22X1 _09104_ (
    .A(_02962_),
    .B(_02385_),
    .C(_02394_),
    .D(_02395_),
    .Y(_02145_)
  );
  NOR2X1 _09105_ (
    .A(execution_unit_0.register_file_0.r9_4_ ),
    .B(_02386_),
    .Y(_02396_)
  );
  OAI21X1 _09106_ (
    .A(_03122_),
    .B(_02387_),
    .C(_02385_),
    .Y(_02397_)
  );
  OAI22X1 _09107_ (
    .A(_02965_),
    .B(_02385_),
    .C(_02396_),
    .D(_02397_),
    .Y(_02146_)
  );
  NOR2X1 _09108_ (
    .A(execution_unit_0.register_file_0.r9_5_ ),
    .B(_02386_),
    .Y(_02398_)
  );
  OAI21X1 _09109_ (
    .A(_03140_),
    .B(_02387_),
    .C(_02385_),
    .Y(_02399_)
  );
  OAI22X1 _09110_ (
    .A(_02966_),
    .B(_02385_),
    .C(_02398_),
    .D(_02399_),
    .Y(_02147_)
  );
  AOI21X1 _09111_ (
    .A(_03157_),
    .B(_02386_),
    .C(_02384_),
    .Y(_02400_)
  );
  OAI21X1 _09112_ (
    .A(execution_unit_0.register_file_0.r9_6_ ),
    .B(_02386_),
    .C(_02400_),
    .Y(_02401_)
  );
  OAI21X1 _09113_ (
    .A(_02967_),
    .B(_02385_),
    .C(_02401_),
    .Y(_02148_)
  );
  NOR2X1 _09114_ (
    .A(execution_unit_0.register_file_0.r9_7_ ),
    .B(_02386_),
    .Y(_02402_)
  );
  OAI21X1 _09115_ (
    .A(_03177_),
    .B(_02387_),
    .C(_02385_),
    .Y(_02403_)
  );
  OAI22X1 _09116_ (
    .A(_02968_),
    .B(_02385_),
    .C(_02402_),
    .D(_02403_),
    .Y(_02149_)
  );
  OAI21X1 _09117_ (
    .A(_03195_),
    .B(_02387_),
    .C(_02385_),
    .Y(_02404_)
  );
  INVX1 _09118_ (
    .A(_02404_),
    .Y(_02405_)
  );
  OAI21X1 _09119_ (
    .A(execution_unit_0.register_file_0.r9_8_ ),
    .B(_02386_),
    .C(_02405_),
    .Y(_02406_)
  );
  OAI21X1 _09120_ (
    .A(_02982_),
    .B(_02385_),
    .C(_02406_),
    .Y(_02150_)
  );
  OAI21X1 _09121_ (
    .A(_03212_),
    .B(_02387_),
    .C(_02385_),
    .Y(_02407_)
  );
  INVX1 _09122_ (
    .A(_02407_),
    .Y(_02408_)
  );
  OAI21X1 _09123_ (
    .A(execution_unit_0.register_file_0.r9_9_ ),
    .B(_02386_),
    .C(_02408_),
    .Y(_02409_)
  );
  OAI21X1 _09124_ (
    .A(_02983_),
    .B(_02385_),
    .C(_02409_),
    .Y(_02151_)
  );
  AOI21X1 _09125_ (
    .A(_03231_),
    .B(_02386_),
    .C(_02384_),
    .Y(_02410_)
  );
  OAI21X1 _09126_ (
    .A(execution_unit_0.register_file_0.r9_10_ ),
    .B(_02386_),
    .C(_02410_),
    .Y(_02411_)
  );
  OAI21X1 _09127_ (
    .A(_02984_),
    .B(_02385_),
    .C(_02411_),
    .Y(_02137_)
  );
  OAI21X1 _09128_ (
    .A(execution_unit_0.register_file_0.r9_11_ ),
    .B(_02386_),
    .C(_02385_),
    .Y(_02412_)
  );
  INVX1 _09129_ (
    .A(_02412_),
    .Y(_02413_)
  );
  OAI21X1 _09130_ (
    .A(_03249_),
    .B(_02387_),
    .C(_02413_),
    .Y(_02414_)
  );
  OAI21X1 _09131_ (
    .A(_02985_),
    .B(_02385_),
    .C(_02414_),
    .Y(_02138_)
  );
  OAI21X1 _09132_ (
    .A(execution_unit_0.register_file_0.r9_12_ ),
    .B(_02386_),
    .C(_02385_),
    .Y(_02415_)
  );
  INVX1 _09133_ (
    .A(_02415_),
    .Y(_02416_)
  );
  OAI21X1 _09134_ (
    .A(_03267_),
    .B(_02387_),
    .C(_02416_),
    .Y(_02417_)
  );
  OAI21X1 _09135_ (
    .A(_02986_),
    .B(_02385_),
    .C(_02417_),
    .Y(_02139_)
  );
  OAI21X1 _09136_ (
    .A(execution_unit_0.register_file_0.r9_13_ ),
    .B(_02386_),
    .C(_02385_),
    .Y(_02418_)
  );
  INVX1 _09137_ (
    .A(_02418_),
    .Y(_02419_)
  );
  OAI21X1 _09138_ (
    .A(_03285_),
    .B(_02387_),
    .C(_02419_),
    .Y(_02420_)
  );
  OAI21X1 _09139_ (
    .A(_02987_),
    .B(_02385_),
    .C(_02420_),
    .Y(_02140_)
  );
  OAI21X1 _09140_ (
    .A(execution_unit_0.register_file_0.r9_14_ ),
    .B(_02386_),
    .C(_02385_),
    .Y(_02421_)
  );
  INVX1 _09141_ (
    .A(_02421_),
    .Y(_02422_)
  );
  OAI21X1 _09142_ (
    .A(_03303_),
    .B(_02387_),
    .C(_02422_),
    .Y(_02423_)
  );
  OAI21X1 _09143_ (
    .A(_02988_),
    .B(_02385_),
    .C(_02423_),
    .Y(_02141_)
  );
  OAI21X1 _09144_ (
    .A(execution_unit_0.register_file_0.r9_15_ ),
    .B(_02386_),
    .C(_02385_),
    .Y(_02424_)
  );
  INVX1 _09145_ (
    .A(_02424_),
    .Y(_02425_)
  );
  OAI21X1 _09146_ (
    .A(_02165_),
    .B(_02387_),
    .C(_02425_),
    .Y(_02426_)
  );
  OAI21X1 _09147_ (
    .A(_02989_),
    .B(_02385_),
    .C(_02426_),
    .Y(_02142_)
  );
  AND2X1 _09148_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_8_ ),
    .Y(_02427_)
  );
  NAND2X1 _09149_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_8_ ),
    .Y(_02428_)
  );
  AND2X1 _09150_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03022_),
    .Y(_02429_)
  );
  NAND2X1 _09151_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03022_),
    .Y(_02430_)
  );
  AOI21X1 _09152_ (
    .A(_03037_),
    .B(_02429_),
    .C(_02427_),
    .Y(_02431_)
  );
  OAI21X1 _09153_ (
    .A(execution_unit_0.register_file_0.r8_0_ ),
    .B(_02429_),
    .C(_02431_),
    .Y(_02432_)
  );
  OAI21X1 _09154_ (
    .A(_02955_),
    .B(_02428_),
    .C(_02432_),
    .Y(_02120_)
  );
  NOR2X1 _09155_ (
    .A(execution_unit_0.register_file_0.r8_1_ ),
    .B(_02429_),
    .Y(_02433_)
  );
  OAI21X1 _09156_ (
    .A(_03062_),
    .B(_02430_),
    .C(_02428_),
    .Y(_02434_)
  );
  OAI22X1 _09157_ (
    .A(_02956_),
    .B(_02428_),
    .C(_02433_),
    .D(_02434_),
    .Y(_02127_)
  );
  AOI21X1 _09158_ (
    .A(_03083_),
    .B(_02429_),
    .C(_02427_),
    .Y(_02435_)
  );
  OAI21X1 _09159_ (
    .A(execution_unit_0.register_file_0.r8_2_ ),
    .B(_02429_),
    .C(_02435_),
    .Y(_02436_)
  );
  OAI21X1 _09160_ (
    .A(_02959_),
    .B(_02428_),
    .C(_02436_),
    .Y(_02128_)
  );
  NOR2X1 _09161_ (
    .A(execution_unit_0.register_file_0.r8_3_ ),
    .B(_02429_),
    .Y(_02437_)
  );
  OAI21X1 _09162_ (
    .A(_03104_),
    .B(_02430_),
    .C(_02428_),
    .Y(_02438_)
  );
  OAI22X1 _09163_ (
    .A(_02962_),
    .B(_02428_),
    .C(_02437_),
    .D(_02438_),
    .Y(_02129_)
  );
  NOR2X1 _09164_ (
    .A(execution_unit_0.register_file_0.r8_4_ ),
    .B(_02429_),
    .Y(_02439_)
  );
  OAI21X1 _09165_ (
    .A(_03122_),
    .B(_02430_),
    .C(_02428_),
    .Y(_02440_)
  );
  OAI22X1 _09166_ (
    .A(_02965_),
    .B(_02428_),
    .C(_02439_),
    .D(_02440_),
    .Y(_02130_)
  );
  NOR2X1 _09167_ (
    .A(execution_unit_0.register_file_0.r8_5_ ),
    .B(_02429_),
    .Y(_02441_)
  );
  OAI21X1 _09168_ (
    .A(_03140_),
    .B(_02430_),
    .C(_02428_),
    .Y(_02442_)
  );
  OAI22X1 _09169_ (
    .A(_02966_),
    .B(_02428_),
    .C(_02441_),
    .D(_02442_),
    .Y(_02131_)
  );
  AOI21X1 _09170_ (
    .A(_03157_),
    .B(_02429_),
    .C(_02427_),
    .Y(_02443_)
  );
  OAI21X1 _09171_ (
    .A(execution_unit_0.register_file_0.r8_6_ ),
    .B(_02429_),
    .C(_02443_),
    .Y(_02444_)
  );
  OAI21X1 _09172_ (
    .A(_02967_),
    .B(_02428_),
    .C(_02444_),
    .Y(_02132_)
  );
  NOR2X1 _09173_ (
    .A(execution_unit_0.register_file_0.r8_7_ ),
    .B(_02429_),
    .Y(_02445_)
  );
  OAI21X1 _09174_ (
    .A(_03177_),
    .B(_02430_),
    .C(_02428_),
    .Y(_02446_)
  );
  OAI22X1 _09175_ (
    .A(_02968_),
    .B(_02428_),
    .C(_02445_),
    .D(_02446_),
    .Y(_02133_)
  );
  OAI21X1 _09176_ (
    .A(_03195_),
    .B(_02430_),
    .C(_02428_),
    .Y(_02447_)
  );
  INVX1 _09177_ (
    .A(_02447_),
    .Y(_02448_)
  );
  OAI21X1 _09178_ (
    .A(execution_unit_0.register_file_0.r8_8_ ),
    .B(_02429_),
    .C(_02448_),
    .Y(_02449_)
  );
  OAI21X1 _09179_ (
    .A(_02982_),
    .B(_02428_),
    .C(_02449_),
    .Y(_02134_)
  );
  OAI21X1 _09180_ (
    .A(_03212_),
    .B(_02430_),
    .C(_02428_),
    .Y(_02450_)
  );
  INVX1 _09181_ (
    .A(_02450_),
    .Y(_02451_)
  );
  OAI21X1 _09182_ (
    .A(execution_unit_0.register_file_0.r8_9_ ),
    .B(_02429_),
    .C(_02451_),
    .Y(_02452_)
  );
  OAI21X1 _09183_ (
    .A(_02983_),
    .B(_02428_),
    .C(_02452_),
    .Y(_02135_)
  );
  AOI21X1 _09184_ (
    .A(_03231_),
    .B(_02429_),
    .C(_02427_),
    .Y(_02453_)
  );
  OAI21X1 _09185_ (
    .A(execution_unit_0.register_file_0.r8_10_ ),
    .B(_02429_),
    .C(_02453_),
    .Y(_02454_)
  );
  OAI21X1 _09186_ (
    .A(_02984_),
    .B(_02428_),
    .C(_02454_),
    .Y(_02121_)
  );
  OAI21X1 _09187_ (
    .A(execution_unit_0.register_file_0.r8_11_ ),
    .B(_02429_),
    .C(_02428_),
    .Y(_02455_)
  );
  INVX1 _09188_ (
    .A(_02455_),
    .Y(_02456_)
  );
  OAI21X1 _09189_ (
    .A(_03249_),
    .B(_02430_),
    .C(_02456_),
    .Y(_02457_)
  );
  OAI21X1 _09190_ (
    .A(_02985_),
    .B(_02428_),
    .C(_02457_),
    .Y(_02122_)
  );
  OAI21X1 _09191_ (
    .A(execution_unit_0.register_file_0.r8_12_ ),
    .B(_02429_),
    .C(_02428_),
    .Y(_02458_)
  );
  INVX1 _09192_ (
    .A(_02458_),
    .Y(_02459_)
  );
  OAI21X1 _09193_ (
    .A(_03267_),
    .B(_02430_),
    .C(_02459_),
    .Y(_02460_)
  );
  OAI21X1 _09194_ (
    .A(_02986_),
    .B(_02428_),
    .C(_02460_),
    .Y(_02123_)
  );
  OAI21X1 _09195_ (
    .A(execution_unit_0.register_file_0.r8_13_ ),
    .B(_02429_),
    .C(_02428_),
    .Y(_02461_)
  );
  INVX1 _09196_ (
    .A(_02461_),
    .Y(_02462_)
  );
  OAI21X1 _09197_ (
    .A(_03285_),
    .B(_02430_),
    .C(_02462_),
    .Y(_02463_)
  );
  OAI21X1 _09198_ (
    .A(_02987_),
    .B(_02428_),
    .C(_02463_),
    .Y(_02124_)
  );
  OAI21X1 _09199_ (
    .A(execution_unit_0.register_file_0.r8_14_ ),
    .B(_02429_),
    .C(_02428_),
    .Y(_02464_)
  );
  INVX1 _09200_ (
    .A(_02464_),
    .Y(_02465_)
  );
  OAI21X1 _09201_ (
    .A(_03303_),
    .B(_02430_),
    .C(_02465_),
    .Y(_02466_)
  );
  OAI21X1 _09202_ (
    .A(_02988_),
    .B(_02428_),
    .C(_02466_),
    .Y(_02125_)
  );
  OAI21X1 _09203_ (
    .A(execution_unit_0.register_file_0.r8_15_ ),
    .B(_02429_),
    .C(_02428_),
    .Y(_02467_)
  );
  INVX1 _09204_ (
    .A(_02467_),
    .Y(_02468_)
  );
  OAI21X1 _09205_ (
    .A(_02165_),
    .B(_02430_),
    .C(_02468_),
    .Y(_02469_)
  );
  OAI21X1 _09206_ (
    .A(_02989_),
    .B(_02428_),
    .C(_02469_),
    .Y(_02126_)
  );
  AND2X1 _09207_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_7_ ),
    .Y(_02470_)
  );
  NAND2X1 _09208_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_7_ ),
    .Y(_02471_)
  );
  AND2X1 _09209_ (
    .A(execution_unit_0.reg_incr ),
    .B(_02995_),
    .Y(_02472_)
  );
  NAND2X1 _09210_ (
    .A(execution_unit_0.reg_incr ),
    .B(_02995_),
    .Y(_02473_)
  );
  AOI21X1 _09211_ (
    .A(_03037_),
    .B(_02472_),
    .C(_02470_),
    .Y(_02474_)
  );
  OAI21X1 _09212_ (
    .A(execution_unit_0.register_file_0.r7_0_ ),
    .B(_02472_),
    .C(_02474_),
    .Y(_02475_)
  );
  OAI21X1 _09213_ (
    .A(_02955_),
    .B(_02471_),
    .C(_02475_),
    .Y(_02104_)
  );
  NOR2X1 _09214_ (
    .A(execution_unit_0.register_file_0.r7_1_ ),
    .B(_02472_),
    .Y(_02476_)
  );
  OAI21X1 _09215_ (
    .A(_03062_),
    .B(_02473_),
    .C(_02471_),
    .Y(_02477_)
  );
  OAI22X1 _09216_ (
    .A(_02956_),
    .B(_02471_),
    .C(_02476_),
    .D(_02477_),
    .Y(_02111_)
  );
  AOI21X1 _09217_ (
    .A(_03083_),
    .B(_02472_),
    .C(_02470_),
    .Y(_02478_)
  );
  OAI21X1 _09218_ (
    .A(execution_unit_0.register_file_0.r7_2_ ),
    .B(_02472_),
    .C(_02478_),
    .Y(_02479_)
  );
  OAI21X1 _09219_ (
    .A(_02959_),
    .B(_02471_),
    .C(_02479_),
    .Y(_02112_)
  );
  NOR2X1 _09220_ (
    .A(execution_unit_0.register_file_0.r7_3_ ),
    .B(_02472_),
    .Y(_02480_)
  );
  OAI21X1 _09221_ (
    .A(_03104_),
    .B(_02473_),
    .C(_02471_),
    .Y(_02481_)
  );
  OAI22X1 _09222_ (
    .A(_02962_),
    .B(_02471_),
    .C(_02480_),
    .D(_02481_),
    .Y(_02113_)
  );
  NOR2X1 _09223_ (
    .A(execution_unit_0.register_file_0.r7_4_ ),
    .B(_02472_),
    .Y(_02482_)
  );
  OAI21X1 _09224_ (
    .A(_03122_),
    .B(_02473_),
    .C(_02471_),
    .Y(_02483_)
  );
  OAI22X1 _09225_ (
    .A(_02965_),
    .B(_02471_),
    .C(_02482_),
    .D(_02483_),
    .Y(_02114_)
  );
  NOR2X1 _09226_ (
    .A(execution_unit_0.register_file_0.r7_5_ ),
    .B(_02472_),
    .Y(_02484_)
  );
  OAI21X1 _09227_ (
    .A(_03140_),
    .B(_02473_),
    .C(_02471_),
    .Y(_02485_)
  );
  OAI22X1 _09228_ (
    .A(_02966_),
    .B(_02471_),
    .C(_02484_),
    .D(_02485_),
    .Y(_02115_)
  );
  AOI21X1 _09229_ (
    .A(_03157_),
    .B(_02472_),
    .C(_02470_),
    .Y(_02486_)
  );
  OAI21X1 _09230_ (
    .A(execution_unit_0.register_file_0.r7_6_ ),
    .B(_02472_),
    .C(_02486_),
    .Y(_02487_)
  );
  OAI21X1 _09231_ (
    .A(_02967_),
    .B(_02471_),
    .C(_02487_),
    .Y(_02116_)
  );
  NOR2X1 _09232_ (
    .A(execution_unit_0.register_file_0.r7_7_ ),
    .B(_02472_),
    .Y(_02488_)
  );
  OAI21X1 _09233_ (
    .A(_03177_),
    .B(_02473_),
    .C(_02471_),
    .Y(_02489_)
  );
  OAI22X1 _09234_ (
    .A(_02968_),
    .B(_02471_),
    .C(_02488_),
    .D(_02489_),
    .Y(_02117_)
  );
  OAI21X1 _09235_ (
    .A(_03195_),
    .B(_02473_),
    .C(_02471_),
    .Y(_02490_)
  );
  INVX1 _09236_ (
    .A(_02490_),
    .Y(_02491_)
  );
  OAI21X1 _09237_ (
    .A(execution_unit_0.register_file_0.r7_8_ ),
    .B(_02472_),
    .C(_02491_),
    .Y(_02492_)
  );
  OAI21X1 _09238_ (
    .A(_02982_),
    .B(_02471_),
    .C(_02492_),
    .Y(_02118_)
  );
  OAI21X1 _09239_ (
    .A(_03212_),
    .B(_02473_),
    .C(_02471_),
    .Y(_02493_)
  );
  INVX1 _09240_ (
    .A(_02493_),
    .Y(_02494_)
  );
  OAI21X1 _09241_ (
    .A(execution_unit_0.register_file_0.r7_9_ ),
    .B(_02472_),
    .C(_02494_),
    .Y(_02495_)
  );
  OAI21X1 _09242_ (
    .A(_02983_),
    .B(_02471_),
    .C(_02495_),
    .Y(_02119_)
  );
  AOI21X1 _09243_ (
    .A(_03231_),
    .B(_02472_),
    .C(_02470_),
    .Y(_02496_)
  );
  OAI21X1 _09244_ (
    .A(execution_unit_0.register_file_0.r7_10_ ),
    .B(_02472_),
    .C(_02496_),
    .Y(_02497_)
  );
  OAI21X1 _09245_ (
    .A(_02984_),
    .B(_02471_),
    .C(_02497_),
    .Y(_02105_)
  );
  OAI21X1 _09246_ (
    .A(execution_unit_0.register_file_0.r7_11_ ),
    .B(_02472_),
    .C(_02471_),
    .Y(_02498_)
  );
  INVX1 _09247_ (
    .A(_02498_),
    .Y(_02499_)
  );
  OAI21X1 _09248_ (
    .A(_03249_),
    .B(_02473_),
    .C(_02499_),
    .Y(_02500_)
  );
  OAI21X1 _09249_ (
    .A(_02985_),
    .B(_02471_),
    .C(_02500_),
    .Y(_02106_)
  );
  OAI21X1 _09250_ (
    .A(execution_unit_0.register_file_0.r7_12_ ),
    .B(_02472_),
    .C(_02471_),
    .Y(_02501_)
  );
  INVX1 _09251_ (
    .A(_02501_),
    .Y(_02502_)
  );
  OAI21X1 _09252_ (
    .A(_03267_),
    .B(_02473_),
    .C(_02502_),
    .Y(_02503_)
  );
  OAI21X1 _09253_ (
    .A(_02986_),
    .B(_02471_),
    .C(_02503_),
    .Y(_02107_)
  );
  OAI21X1 _09254_ (
    .A(execution_unit_0.register_file_0.r7_13_ ),
    .B(_02472_),
    .C(_02471_),
    .Y(_02504_)
  );
  INVX1 _09255_ (
    .A(_02504_),
    .Y(_02505_)
  );
  OAI21X1 _09256_ (
    .A(_03285_),
    .B(_02473_),
    .C(_02505_),
    .Y(_02506_)
  );
  OAI21X1 _09257_ (
    .A(_02987_),
    .B(_02471_),
    .C(_02506_),
    .Y(_02108_)
  );
  OAI21X1 _09258_ (
    .A(execution_unit_0.register_file_0.r7_14_ ),
    .B(_02472_),
    .C(_02471_),
    .Y(_02507_)
  );
  INVX1 _09259_ (
    .A(_02507_),
    .Y(_02508_)
  );
  OAI21X1 _09260_ (
    .A(_03303_),
    .B(_02473_),
    .C(_02508_),
    .Y(_02509_)
  );
  OAI21X1 _09261_ (
    .A(_02988_),
    .B(_02471_),
    .C(_02509_),
    .Y(_02109_)
  );
  OAI21X1 _09262_ (
    .A(execution_unit_0.register_file_0.r7_15_ ),
    .B(_02472_),
    .C(_02471_),
    .Y(_02510_)
  );
  INVX1 _09263_ (
    .A(_02510_),
    .Y(_02511_)
  );
  OAI21X1 _09264_ (
    .A(_02165_),
    .B(_02473_),
    .C(_02511_),
    .Y(_02512_)
  );
  OAI21X1 _09265_ (
    .A(_02989_),
    .B(_02471_),
    .C(_02512_),
    .Y(_02110_)
  );
  AND2X1 _09266_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_6_ ),
    .Y(_02513_)
  );
  NAND2X1 _09267_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_6_ ),
    .Y(_02514_)
  );
  AND2X1 _09268_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03013_),
    .Y(_02515_)
  );
  NAND2X1 _09269_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03013_),
    .Y(_02516_)
  );
  AOI21X1 _09270_ (
    .A(_03037_),
    .B(_02515_),
    .C(_02513_),
    .Y(_02517_)
  );
  OAI21X1 _09271_ (
    .A(execution_unit_0.register_file_0.r6_0_ ),
    .B(_02515_),
    .C(_02517_),
    .Y(_02518_)
  );
  OAI21X1 _09272_ (
    .A(_02955_),
    .B(_02514_),
    .C(_02518_),
    .Y(_02088_)
  );
  NOR2X1 _09273_ (
    .A(execution_unit_0.register_file_0.r6_1_ ),
    .B(_02515_),
    .Y(_02519_)
  );
  OAI21X1 _09274_ (
    .A(_03062_),
    .B(_02516_),
    .C(_02514_),
    .Y(_02520_)
  );
  OAI22X1 _09275_ (
    .A(_02956_),
    .B(_02514_),
    .C(_02519_),
    .D(_02520_),
    .Y(_02095_)
  );
  AOI21X1 _09276_ (
    .A(_03083_),
    .B(_02515_),
    .C(_02513_),
    .Y(_02521_)
  );
  OAI21X1 _09277_ (
    .A(execution_unit_0.register_file_0.r6_2_ ),
    .B(_02515_),
    .C(_02521_),
    .Y(_02522_)
  );
  OAI21X1 _09278_ (
    .A(_02959_),
    .B(_02514_),
    .C(_02522_),
    .Y(_02096_)
  );
  NOR2X1 _09279_ (
    .A(execution_unit_0.register_file_0.r6_3_ ),
    .B(_02515_),
    .Y(_02523_)
  );
  OAI21X1 _09280_ (
    .A(_03104_),
    .B(_02516_),
    .C(_02514_),
    .Y(_02524_)
  );
  OAI22X1 _09281_ (
    .A(_02962_),
    .B(_02514_),
    .C(_02523_),
    .D(_02524_),
    .Y(_02097_)
  );
  NOR2X1 _09282_ (
    .A(execution_unit_0.register_file_0.r6_4_ ),
    .B(_02515_),
    .Y(_02525_)
  );
  OAI21X1 _09283_ (
    .A(_03122_),
    .B(_02516_),
    .C(_02514_),
    .Y(_02526_)
  );
  OAI22X1 _09284_ (
    .A(_02965_),
    .B(_02514_),
    .C(_02525_),
    .D(_02526_),
    .Y(_02098_)
  );
  NOR2X1 _09285_ (
    .A(execution_unit_0.register_file_0.r6_5_ ),
    .B(_02515_),
    .Y(_02527_)
  );
  OAI21X1 _09286_ (
    .A(_03140_),
    .B(_02516_),
    .C(_02514_),
    .Y(_02528_)
  );
  OAI22X1 _09287_ (
    .A(_02966_),
    .B(_02514_),
    .C(_02527_),
    .D(_02528_),
    .Y(_02099_)
  );
  AOI21X1 _09288_ (
    .A(_03157_),
    .B(_02515_),
    .C(_02513_),
    .Y(_02529_)
  );
  OAI21X1 _09289_ (
    .A(execution_unit_0.register_file_0.r6_6_ ),
    .B(_02515_),
    .C(_02529_),
    .Y(_02530_)
  );
  OAI21X1 _09290_ (
    .A(_02967_),
    .B(_02514_),
    .C(_02530_),
    .Y(_02100_)
  );
  NOR2X1 _09291_ (
    .A(execution_unit_0.register_file_0.r6_7_ ),
    .B(_02515_),
    .Y(_02531_)
  );
  OAI21X1 _09292_ (
    .A(_03177_),
    .B(_02516_),
    .C(_02514_),
    .Y(_02532_)
  );
  OAI22X1 _09293_ (
    .A(_02968_),
    .B(_02514_),
    .C(_02531_),
    .D(_02532_),
    .Y(_02101_)
  );
  OAI21X1 _09294_ (
    .A(_03195_),
    .B(_02516_),
    .C(_02514_),
    .Y(_02533_)
  );
  INVX1 _09295_ (
    .A(_02533_),
    .Y(_02534_)
  );
  OAI21X1 _09296_ (
    .A(execution_unit_0.register_file_0.r6_8_ ),
    .B(_02515_),
    .C(_02534_),
    .Y(_02535_)
  );
  OAI21X1 _09297_ (
    .A(_02982_),
    .B(_02514_),
    .C(_02535_),
    .Y(_02102_)
  );
  OAI21X1 _09298_ (
    .A(_03212_),
    .B(_02516_),
    .C(_02514_),
    .Y(_02536_)
  );
  INVX1 _09299_ (
    .A(_02536_),
    .Y(_02537_)
  );
  OAI21X1 _09300_ (
    .A(execution_unit_0.register_file_0.r6_9_ ),
    .B(_02515_),
    .C(_02537_),
    .Y(_02538_)
  );
  OAI21X1 _09301_ (
    .A(_02983_),
    .B(_02514_),
    .C(_02538_),
    .Y(_02103_)
  );
  AOI21X1 _09302_ (
    .A(_03231_),
    .B(_02515_),
    .C(_02513_),
    .Y(_02539_)
  );
  OAI21X1 _09303_ (
    .A(execution_unit_0.register_file_0.r6_10_ ),
    .B(_02515_),
    .C(_02539_),
    .Y(_02540_)
  );
  OAI21X1 _09304_ (
    .A(_02984_),
    .B(_02514_),
    .C(_02540_),
    .Y(_02089_)
  );
  OAI21X1 _09305_ (
    .A(execution_unit_0.register_file_0.r6_11_ ),
    .B(_02515_),
    .C(_02514_),
    .Y(_02541_)
  );
  INVX1 _09306_ (
    .A(_02541_),
    .Y(_02542_)
  );
  OAI21X1 _09307_ (
    .A(_03249_),
    .B(_02516_),
    .C(_02542_),
    .Y(_02543_)
  );
  OAI21X1 _09308_ (
    .A(_02985_),
    .B(_02514_),
    .C(_02543_),
    .Y(_02090_)
  );
  OAI21X1 _09309_ (
    .A(execution_unit_0.register_file_0.r6_12_ ),
    .B(_02515_),
    .C(_02514_),
    .Y(_02544_)
  );
  INVX1 _09310_ (
    .A(_02544_),
    .Y(_02545_)
  );
  OAI21X1 _09311_ (
    .A(_03267_),
    .B(_02516_),
    .C(_02545_),
    .Y(_02546_)
  );
  OAI21X1 _09312_ (
    .A(_02986_),
    .B(_02514_),
    .C(_02546_),
    .Y(_02091_)
  );
  OAI21X1 _09313_ (
    .A(execution_unit_0.register_file_0.r6_13_ ),
    .B(_02515_),
    .C(_02514_),
    .Y(_02547_)
  );
  INVX1 _09314_ (
    .A(_02547_),
    .Y(_02548_)
  );
  OAI21X1 _09315_ (
    .A(_03285_),
    .B(_02516_),
    .C(_02548_),
    .Y(_02549_)
  );
  OAI21X1 _09316_ (
    .A(_02987_),
    .B(_02514_),
    .C(_02549_),
    .Y(_02092_)
  );
  OAI21X1 _09317_ (
    .A(execution_unit_0.register_file_0.r6_14_ ),
    .B(_02515_),
    .C(_02514_),
    .Y(_02550_)
  );
  INVX1 _09318_ (
    .A(_02550_),
    .Y(_02551_)
  );
  OAI21X1 _09319_ (
    .A(_03303_),
    .B(_02516_),
    .C(_02551_),
    .Y(_02552_)
  );
  OAI21X1 _09320_ (
    .A(_02988_),
    .B(_02514_),
    .C(_02552_),
    .Y(_02093_)
  );
  OAI21X1 _09321_ (
    .A(execution_unit_0.register_file_0.r6_15_ ),
    .B(_02515_),
    .C(_02514_),
    .Y(_02553_)
  );
  INVX1 _09322_ (
    .A(_02553_),
    .Y(_02554_)
  );
  OAI21X1 _09323_ (
    .A(_02165_),
    .B(_02516_),
    .C(_02554_),
    .Y(_02555_)
  );
  OAI21X1 _09324_ (
    .A(_02989_),
    .B(_02514_),
    .C(_02555_),
    .Y(_02094_)
  );
  AND2X1 _09325_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_5_ ),
    .Y(_02556_)
  );
  NAND2X1 _09326_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_5_ ),
    .Y(_02557_)
  );
  AND2X1 _09327_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03004_),
    .Y(_02558_)
  );
  NAND2X1 _09328_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03004_),
    .Y(_02559_)
  );
  AOI21X1 _09329_ (
    .A(_03037_),
    .B(_02558_),
    .C(_02556_),
    .Y(_02560_)
  );
  OAI21X1 _09330_ (
    .A(execution_unit_0.register_file_0.r5_0_ ),
    .B(_02558_),
    .C(_02560_),
    .Y(_02561_)
  );
  OAI21X1 _09331_ (
    .A(_02955_),
    .B(_02557_),
    .C(_02561_),
    .Y(_02072_)
  );
  NOR2X1 _09332_ (
    .A(execution_unit_0.register_file_0.r5_1_ ),
    .B(_02558_),
    .Y(_02562_)
  );
  OAI21X1 _09333_ (
    .A(_03062_),
    .B(_02559_),
    .C(_02557_),
    .Y(_02563_)
  );
  OAI22X1 _09334_ (
    .A(_02956_),
    .B(_02557_),
    .C(_02562_),
    .D(_02563_),
    .Y(_02079_)
  );
  AOI21X1 _09335_ (
    .A(_03083_),
    .B(_02558_),
    .C(_02556_),
    .Y(_02564_)
  );
  OAI21X1 _09336_ (
    .A(execution_unit_0.register_file_0.r5_2_ ),
    .B(_02558_),
    .C(_02564_),
    .Y(_02565_)
  );
  OAI21X1 _09337_ (
    .A(_02959_),
    .B(_02557_),
    .C(_02565_),
    .Y(_02080_)
  );
  NOR2X1 _09338_ (
    .A(execution_unit_0.register_file_0.r5_3_ ),
    .B(_02558_),
    .Y(_02566_)
  );
  OAI21X1 _09339_ (
    .A(_03104_),
    .B(_02559_),
    .C(_02557_),
    .Y(_02567_)
  );
  OAI22X1 _09340_ (
    .A(_02962_),
    .B(_02557_),
    .C(_02566_),
    .D(_02567_),
    .Y(_02081_)
  );
  NOR2X1 _09341_ (
    .A(execution_unit_0.register_file_0.r5_4_ ),
    .B(_02558_),
    .Y(_02568_)
  );
  OAI21X1 _09342_ (
    .A(_03122_),
    .B(_02559_),
    .C(_02557_),
    .Y(_02569_)
  );
  OAI22X1 _09343_ (
    .A(_02965_),
    .B(_02557_),
    .C(_02568_),
    .D(_02569_),
    .Y(_02082_)
  );
  NOR2X1 _09344_ (
    .A(execution_unit_0.register_file_0.r5_5_ ),
    .B(_02558_),
    .Y(_02570_)
  );
  OAI21X1 _09345_ (
    .A(_03140_),
    .B(_02559_),
    .C(_02557_),
    .Y(_02571_)
  );
  OAI22X1 _09346_ (
    .A(_02966_),
    .B(_02557_),
    .C(_02570_),
    .D(_02571_),
    .Y(_02083_)
  );
  AOI21X1 _09347_ (
    .A(_03157_),
    .B(_02558_),
    .C(_02556_),
    .Y(_02572_)
  );
  OAI21X1 _09348_ (
    .A(execution_unit_0.register_file_0.r5_6_ ),
    .B(_02558_),
    .C(_02572_),
    .Y(_02573_)
  );
  OAI21X1 _09349_ (
    .A(_02967_),
    .B(_02557_),
    .C(_02573_),
    .Y(_02084_)
  );
  NOR2X1 _09350_ (
    .A(execution_unit_0.register_file_0.r5_7_ ),
    .B(_02558_),
    .Y(_02574_)
  );
  OAI21X1 _09351_ (
    .A(_03177_),
    .B(_02559_),
    .C(_02557_),
    .Y(_02575_)
  );
  OAI22X1 _09352_ (
    .A(_02968_),
    .B(_02557_),
    .C(_02574_),
    .D(_02575_),
    .Y(_02085_)
  );
  OAI21X1 _09353_ (
    .A(_03195_),
    .B(_02559_),
    .C(_02557_),
    .Y(_02576_)
  );
  INVX1 _09354_ (
    .A(_02576_),
    .Y(_02577_)
  );
  OAI21X1 _09355_ (
    .A(execution_unit_0.register_file_0.r5_8_ ),
    .B(_02558_),
    .C(_02577_),
    .Y(_02578_)
  );
  OAI21X1 _09356_ (
    .A(_02982_),
    .B(_02557_),
    .C(_02578_),
    .Y(_02086_)
  );
  OAI21X1 _09357_ (
    .A(_03212_),
    .B(_02559_),
    .C(_02557_),
    .Y(_02579_)
  );
  INVX1 _09358_ (
    .A(_02579_),
    .Y(_02580_)
  );
  OAI21X1 _09359_ (
    .A(execution_unit_0.register_file_0.r5_9_ ),
    .B(_02558_),
    .C(_02580_),
    .Y(_02581_)
  );
  OAI21X1 _09360_ (
    .A(_02983_),
    .B(_02557_),
    .C(_02581_),
    .Y(_02087_)
  );
  AOI21X1 _09361_ (
    .A(_03231_),
    .B(_02558_),
    .C(_02556_),
    .Y(_02582_)
  );
  OAI21X1 _09362_ (
    .A(execution_unit_0.register_file_0.r5_10_ ),
    .B(_02558_),
    .C(_02582_),
    .Y(_02583_)
  );
  OAI21X1 _09363_ (
    .A(_02984_),
    .B(_02557_),
    .C(_02583_),
    .Y(_02073_)
  );
  OAI21X1 _09364_ (
    .A(execution_unit_0.register_file_0.r5_11_ ),
    .B(_02558_),
    .C(_02557_),
    .Y(_02584_)
  );
  INVX1 _09365_ (
    .A(_02584_),
    .Y(_02585_)
  );
  OAI21X1 _09366_ (
    .A(_03249_),
    .B(_02559_),
    .C(_02585_),
    .Y(_02586_)
  );
  OAI21X1 _09367_ (
    .A(_02985_),
    .B(_02557_),
    .C(_02586_),
    .Y(_02074_)
  );
  OAI21X1 _09368_ (
    .A(execution_unit_0.register_file_0.r5_12_ ),
    .B(_02558_),
    .C(_02557_),
    .Y(_02587_)
  );
  INVX1 _09369_ (
    .A(_02587_),
    .Y(_02588_)
  );
  OAI21X1 _09370_ (
    .A(_03267_),
    .B(_02559_),
    .C(_02588_),
    .Y(_02589_)
  );
  OAI21X1 _09371_ (
    .A(_02986_),
    .B(_02557_),
    .C(_02589_),
    .Y(_02075_)
  );
  OAI21X1 _09372_ (
    .A(execution_unit_0.register_file_0.r5_13_ ),
    .B(_02558_),
    .C(_02557_),
    .Y(_02590_)
  );
  INVX1 _09373_ (
    .A(_02590_),
    .Y(_02591_)
  );
  OAI21X1 _09374_ (
    .A(_03285_),
    .B(_02559_),
    .C(_02591_),
    .Y(_02592_)
  );
  OAI21X1 _09375_ (
    .A(_02987_),
    .B(_02557_),
    .C(_02592_),
    .Y(_02076_)
  );
  OAI21X1 _09376_ (
    .A(execution_unit_0.register_file_0.r5_14_ ),
    .B(_02558_),
    .C(_02557_),
    .Y(_02593_)
  );
  INVX1 _09377_ (
    .A(_02593_),
    .Y(_02594_)
  );
  OAI21X1 _09378_ (
    .A(_03303_),
    .B(_02559_),
    .C(_02594_),
    .Y(_02595_)
  );
  OAI21X1 _09379_ (
    .A(_02988_),
    .B(_02557_),
    .C(_02595_),
    .Y(_02077_)
  );
  OAI21X1 _09380_ (
    .A(execution_unit_0.register_file_0.r5_15_ ),
    .B(_02558_),
    .C(_02557_),
    .Y(_02596_)
  );
  INVX1 _09381_ (
    .A(_02596_),
    .Y(_02597_)
  );
  OAI21X1 _09382_ (
    .A(_02165_),
    .B(_02559_),
    .C(_02597_),
    .Y(_02598_)
  );
  OAI21X1 _09383_ (
    .A(_02989_),
    .B(_02557_),
    .C(_02598_),
    .Y(_02078_)
  );
  NAND2X1 _09384_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_3_ ),
    .Y(_02599_)
  );
  NAND2X1 _09385_ (
    .A(execution_unit_0.register_file_0.r3_0_ ),
    .B(_02599_),
    .Y(_02600_)
  );
  OAI21X1 _09386_ (
    .A(_02955_),
    .B(_02599_),
    .C(_02600_),
    .Y(_02040_)
  );
  NAND2X1 _09387_ (
    .A(execution_unit_0.register_file_0.r3_1_ ),
    .B(_02599_),
    .Y(_02601_)
  );
  OAI21X1 _09388_ (
    .A(_02956_),
    .B(_02599_),
    .C(_02601_),
    .Y(_02047_)
  );
  NAND2X1 _09389_ (
    .A(execution_unit_0.register_file_0.r3_2_ ),
    .B(_02599_),
    .Y(_02602_)
  );
  OAI21X1 _09390_ (
    .A(_02959_),
    .B(_02599_),
    .C(_02602_),
    .Y(_02048_)
  );
  NAND2X1 _09391_ (
    .A(execution_unit_0.register_file_0.r3_3_ ),
    .B(_02599_),
    .Y(_02603_)
  );
  OAI21X1 _09392_ (
    .A(_02962_),
    .B(_02599_),
    .C(_02603_),
    .Y(_02049_)
  );
  NAND2X1 _09393_ (
    .A(execution_unit_0.register_file_0.r3_4_ ),
    .B(_02599_),
    .Y(_02604_)
  );
  OAI21X1 _09394_ (
    .A(_02965_),
    .B(_02599_),
    .C(_02604_),
    .Y(_02050_)
  );
  NAND2X1 _09395_ (
    .A(execution_unit_0.register_file_0.r3_5_ ),
    .B(_02599_),
    .Y(_02605_)
  );
  OAI21X1 _09396_ (
    .A(_02966_),
    .B(_02599_),
    .C(_02605_),
    .Y(_02051_)
  );
  NAND2X1 _09397_ (
    .A(execution_unit_0.register_file_0.r3_6_ ),
    .B(_02599_),
    .Y(_02606_)
  );
  OAI21X1 _09398_ (
    .A(_02967_),
    .B(_02599_),
    .C(_02606_),
    .Y(_02052_)
  );
  NAND2X1 _09399_ (
    .A(execution_unit_0.register_file_0.r3_7_ ),
    .B(_02599_),
    .Y(_02607_)
  );
  OAI21X1 _09400_ (
    .A(_02968_),
    .B(_02599_),
    .C(_02607_),
    .Y(_02053_)
  );
  NAND2X1 _09401_ (
    .A(execution_unit_0.register_file_0.r3_8_ ),
    .B(_02599_),
    .Y(_02608_)
  );
  OAI21X1 _09402_ (
    .A(_02982_),
    .B(_02599_),
    .C(_02608_),
    .Y(_02054_)
  );
  NAND2X1 _09403_ (
    .A(execution_unit_0.register_file_0.r3_9_ ),
    .B(_02599_),
    .Y(_02609_)
  );
  OAI21X1 _09404_ (
    .A(_02983_),
    .B(_02599_),
    .C(_02609_),
    .Y(_02055_)
  );
  NAND2X1 _09405_ (
    .A(execution_unit_0.register_file_0.r3_10_ ),
    .B(_02599_),
    .Y(_02610_)
  );
  OAI21X1 _09406_ (
    .A(_02984_),
    .B(_02599_),
    .C(_02610_),
    .Y(_02041_)
  );
  NAND2X1 _09407_ (
    .A(execution_unit_0.register_file_0.r3_11_ ),
    .B(_02599_),
    .Y(_02611_)
  );
  OAI21X1 _09408_ (
    .A(_02985_),
    .B(_02599_),
    .C(_02611_),
    .Y(_02042_)
  );
  NAND2X1 _09409_ (
    .A(execution_unit_0.register_file_0.r3_12_ ),
    .B(_02599_),
    .Y(_02612_)
  );
  OAI21X1 _09410_ (
    .A(_02986_),
    .B(_02599_),
    .C(_02612_),
    .Y(_02043_)
  );
  NAND2X1 _09411_ (
    .A(execution_unit_0.register_file_0.r3_13_ ),
    .B(_02599_),
    .Y(_02613_)
  );
  OAI21X1 _09412_ (
    .A(_02987_),
    .B(_02599_),
    .C(_02613_),
    .Y(_02044_)
  );
  NAND2X1 _09413_ (
    .A(execution_unit_0.register_file_0.r3_14_ ),
    .B(_02599_),
    .Y(_02614_)
  );
  OAI21X1 _09414_ (
    .A(_02988_),
    .B(_02599_),
    .C(_02614_),
    .Y(_02045_)
  );
  NAND2X1 _09415_ (
    .A(execution_unit_0.register_file_0.r3_15_ ),
    .B(_02599_),
    .Y(_02615_)
  );
  OAI21X1 _09416_ (
    .A(_02989_),
    .B(_02599_),
    .C(_02615_),
    .Y(_02046_)
  );
  AND2X1 _09417_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_4_ ),
    .Y(_02616_)
  );
  NAND2X1 _09418_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_4_ ),
    .Y(_02617_)
  );
  AND2X1 _09419_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03007_),
    .Y(_02618_)
  );
  NAND2X1 _09420_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03007_),
    .Y(_02619_)
  );
  AOI21X1 _09421_ (
    .A(_03037_),
    .B(_02618_),
    .C(_02616_),
    .Y(_02620_)
  );
  OAI21X1 _09422_ (
    .A(execution_unit_0.register_file_0.r4_0_ ),
    .B(_02618_),
    .C(_02620_),
    .Y(_02621_)
  );
  OAI21X1 _09423_ (
    .A(_02955_),
    .B(_02617_),
    .C(_02621_),
    .Y(_02056_)
  );
  NOR2X1 _09424_ (
    .A(execution_unit_0.register_file_0.r4_1_ ),
    .B(_02618_),
    .Y(_02622_)
  );
  OAI21X1 _09425_ (
    .A(_03062_),
    .B(_02619_),
    .C(_02617_),
    .Y(_02623_)
  );
  OAI22X1 _09426_ (
    .A(_02956_),
    .B(_02617_),
    .C(_02622_),
    .D(_02623_),
    .Y(_02063_)
  );
  AOI21X1 _09427_ (
    .A(_03083_),
    .B(_02618_),
    .C(_02616_),
    .Y(_02624_)
  );
  OAI21X1 _09428_ (
    .A(execution_unit_0.register_file_0.r4_2_ ),
    .B(_02618_),
    .C(_02624_),
    .Y(_02625_)
  );
  OAI21X1 _09429_ (
    .A(_02959_),
    .B(_02617_),
    .C(_02625_),
    .Y(_02064_)
  );
  NOR2X1 _09430_ (
    .A(execution_unit_0.register_file_0.r4_3_ ),
    .B(_02618_),
    .Y(_02626_)
  );
  OAI21X1 _09431_ (
    .A(_03104_),
    .B(_02619_),
    .C(_02617_),
    .Y(_02627_)
  );
  OAI22X1 _09432_ (
    .A(_02962_),
    .B(_02617_),
    .C(_02626_),
    .D(_02627_),
    .Y(_02065_)
  );
  NOR2X1 _09433_ (
    .A(execution_unit_0.register_file_0.r4_4_ ),
    .B(_02618_),
    .Y(_02628_)
  );
  OAI21X1 _09434_ (
    .A(_03122_),
    .B(_02619_),
    .C(_02617_),
    .Y(_02629_)
  );
  OAI22X1 _09435_ (
    .A(_02965_),
    .B(_02617_),
    .C(_02628_),
    .D(_02629_),
    .Y(_02066_)
  );
  NOR2X1 _09436_ (
    .A(execution_unit_0.register_file_0.r4_5_ ),
    .B(_02618_),
    .Y(_02630_)
  );
  OAI21X1 _09437_ (
    .A(_03140_),
    .B(_02619_),
    .C(_02617_),
    .Y(_02631_)
  );
  OAI22X1 _09438_ (
    .A(_02966_),
    .B(_02617_),
    .C(_02630_),
    .D(_02631_),
    .Y(_02067_)
  );
  AOI21X1 _09439_ (
    .A(_03157_),
    .B(_02618_),
    .C(_02616_),
    .Y(_02632_)
  );
  OAI21X1 _09440_ (
    .A(execution_unit_0.register_file_0.r4_6_ ),
    .B(_02618_),
    .C(_02632_),
    .Y(_02633_)
  );
  OAI21X1 _09441_ (
    .A(_02967_),
    .B(_02617_),
    .C(_02633_),
    .Y(_02068_)
  );
  NOR2X1 _09442_ (
    .A(execution_unit_0.register_file_0.r4_7_ ),
    .B(_02618_),
    .Y(_02634_)
  );
  OAI21X1 _09443_ (
    .A(_03177_),
    .B(_02619_),
    .C(_02617_),
    .Y(_02635_)
  );
  OAI22X1 _09444_ (
    .A(_02968_),
    .B(_02617_),
    .C(_02634_),
    .D(_02635_),
    .Y(_02069_)
  );
  OAI21X1 _09445_ (
    .A(_03195_),
    .B(_02619_),
    .C(_02617_),
    .Y(_02636_)
  );
  INVX1 _09446_ (
    .A(_02636_),
    .Y(_02637_)
  );
  OAI21X1 _09447_ (
    .A(execution_unit_0.register_file_0.r4_8_ ),
    .B(_02618_),
    .C(_02637_),
    .Y(_02638_)
  );
  OAI21X1 _09448_ (
    .A(_02982_),
    .B(_02617_),
    .C(_02638_),
    .Y(_02070_)
  );
  OAI21X1 _09449_ (
    .A(_03212_),
    .B(_02619_),
    .C(_02617_),
    .Y(_02639_)
  );
  INVX1 _09450_ (
    .A(_02639_),
    .Y(_02640_)
  );
  OAI21X1 _09451_ (
    .A(execution_unit_0.register_file_0.r4_9_ ),
    .B(_02618_),
    .C(_02640_),
    .Y(_02641_)
  );
  OAI21X1 _09452_ (
    .A(_02983_),
    .B(_02617_),
    .C(_02641_),
    .Y(_02071_)
  );
  OAI21X1 _09453_ (
    .A(execution_unit_0.register_file_0.r4_10_ ),
    .B(_02618_),
    .C(_02617_),
    .Y(_02642_)
  );
  AOI21X1 _09454_ (
    .A(_03231_),
    .B(_02618_),
    .C(_02642_),
    .Y(_02643_)
  );
  INVX1 _09455_ (
    .A(_02643_),
    .Y(_02644_)
  );
  OAI21X1 _09456_ (
    .A(_02984_),
    .B(_02617_),
    .C(_02644_),
    .Y(_02057_)
  );
  OAI21X1 _09457_ (
    .A(execution_unit_0.register_file_0.r4_11_ ),
    .B(_02618_),
    .C(_02617_),
    .Y(_02645_)
  );
  INVX1 _09458_ (
    .A(_02645_),
    .Y(_02646_)
  );
  OAI21X1 _09459_ (
    .A(_03249_),
    .B(_02619_),
    .C(_02646_),
    .Y(_02647_)
  );
  OAI21X1 _09460_ (
    .A(_02985_),
    .B(_02617_),
    .C(_02647_),
    .Y(_02058_)
  );
  OAI21X1 _09461_ (
    .A(execution_unit_0.register_file_0.r4_12_ ),
    .B(_02618_),
    .C(_02617_),
    .Y(_02648_)
  );
  INVX1 _09462_ (
    .A(_02648_),
    .Y(_02649_)
  );
  OAI21X1 _09463_ (
    .A(_03267_),
    .B(_02619_),
    .C(_02649_),
    .Y(_02650_)
  );
  OAI21X1 _09464_ (
    .A(_02986_),
    .B(_02617_),
    .C(_02650_),
    .Y(_02059_)
  );
  OAI21X1 _09465_ (
    .A(execution_unit_0.register_file_0.r4_13_ ),
    .B(_02618_),
    .C(_02617_),
    .Y(_02651_)
  );
  INVX1 _09466_ (
    .A(_02651_),
    .Y(_02652_)
  );
  OAI21X1 _09467_ (
    .A(_03285_),
    .B(_02619_),
    .C(_02652_),
    .Y(_02653_)
  );
  OAI21X1 _09468_ (
    .A(_02987_),
    .B(_02617_),
    .C(_02653_),
    .Y(_02060_)
  );
  OAI21X1 _09469_ (
    .A(execution_unit_0.register_file_0.r4_14_ ),
    .B(_02618_),
    .C(_02617_),
    .Y(_02654_)
  );
  INVX1 _09470_ (
    .A(_02654_),
    .Y(_02655_)
  );
  OAI21X1 _09471_ (
    .A(_03303_),
    .B(_02619_),
    .C(_02655_),
    .Y(_02656_)
  );
  OAI21X1 _09472_ (
    .A(_02988_),
    .B(_02617_),
    .C(_02656_),
    .Y(_02061_)
  );
  OAI21X1 _09473_ (
    .A(execution_unit_0.register_file_0.r4_15_ ),
    .B(_02618_),
    .C(_02617_),
    .Y(_02657_)
  );
  INVX1 _09474_ (
    .A(_02657_),
    .Y(_02658_)
  );
  OAI21X1 _09475_ (
    .A(_02165_),
    .B(_02619_),
    .C(_02658_),
    .Y(_02659_)
  );
  OAI21X1 _09476_ (
    .A(_02989_),
    .B(_02617_),
    .C(_02659_),
    .Y(_02062_)
  );
  AOI21X1 _09477_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_2_ ),
    .C(execution_unit_0.reg_sr_wr ),
    .Y(_02660_)
  );
  MUX2X1 _09478_ (
    .A(execution_unit_0.alu_0.status_0_ ),
    .B(execution_unit_0.alu_0.alu_out_0_ ),
    .S(_02660_),
    .Y(_02661_)
  );
  OAI21X1 _09479_ (
    .A(execution_unit_0.alu_0.alu_stat_0_ ),
    .B(_02977_),
    .C(_02950_),
    .Y(_02662_)
  );
  AOI21X1 _09480_ (
    .A(_02977_),
    .B(_02661_),
    .C(_02662_),
    .Y(_02032_)
  );
  MUX2X1 _09481_ (
    .A(execution_unit_0.alu_0.status_1_ ),
    .B(execution_unit_0.alu_0.alu_out_1_ ),
    .S(_02660_),
    .Y(_02663_)
  );
  OAI21X1 _09482_ (
    .A(execution_unit_0.alu_0.Z ),
    .B(_02978_),
    .C(_02950_),
    .Y(_02664_)
  );
  AOI21X1 _09483_ (
    .A(_02978_),
    .B(_02663_),
    .C(_02664_),
    .Y(_02033_)
  );
  MUX2X1 _09484_ (
    .A(execution_unit_0.alu_0.status_2_ ),
    .B(execution_unit_0.alu_0.alu_out_2_ ),
    .S(_02660_),
    .Y(_02665_)
  );
  OAI21X1 _09485_ (
    .A(execution_unit_0.alu_0.N ),
    .B(_02979_),
    .C(_02950_),
    .Y(_02666_)
  );
  AOI21X1 _09486_ (
    .A(_02979_),
    .B(_02665_),
    .C(_02666_),
    .Y(_02034_)
  );
  MUX2X1 _09487_ (
    .A(execution_unit_0.gie ),
    .B(execution_unit_0.alu_0.alu_out_3_ ),
    .S(_02660_),
    .Y(_02667_)
  );
  NOR2X1 _09488_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02667_),
    .Y(_02035_)
  );
  OAI21X1 _09489_ (
    .A(_02965_),
    .B(_02660_),
    .C(_02963_),
    .Y(clock_module_0.UNUSED_cpuoff )
  );
  MUX2X1 _09490_ (
    .A(execution_unit_0.register_file_0.r2_4_ ),
    .B(execution_unit_0.alu_0.alu_out_4_ ),
    .S(_02660_),
    .Y(_02668_)
  );
  NOR2X1 _09491_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02668_),
    .Y(_02036_)
  );
  MUX2X1 _09492_ (
    .A(clock_module_0.oscoff ),
    .B(execution_unit_0.alu_0.alu_out_5_ ),
    .S(_02660_),
    .Y(_02669_)
  );
  NOR2X1 _09493_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02669_),
    .Y(_02037_)
  );
  MUX2X1 _09494_ (
    .A(clock_module_0.scg1 ),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .S(_02660_),
    .Y(_02670_)
  );
  NOR2X1 _09495_ (
    .A(execution_unit_0.reg_sr_clr ),
    .B(_02670_),
    .Y(_02038_)
  );
  OAI21X1 _09496_ (
    .A(_02982_),
    .B(_02660_),
    .C(_02980_),
    .Y(_02671_)
  );
  AOI21X1 _09497_ (
    .A(execution_unit_0.alu_0.status_3_ ),
    .B(_02660_),
    .C(_02671_),
    .Y(_02672_)
  );
  OAI21X1 _09498_ (
    .A(execution_unit_0.alu_0.alu_stat_3_ ),
    .B(_02980_),
    .C(_02950_),
    .Y(_02673_)
  );
  NOR2X1 _09499_ (
    .A(_02672_),
    .B(_02673_),
    .Y(_02039_)
  );
  AND2X1 _09500_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03001_),
    .Y(_02674_)
  );
  NAND2X1 _09501_ (
    .A(execution_unit_0.reg_incr ),
    .B(_03001_),
    .Y(_02675_)
  );
  AND2X1 _09502_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_1_ ),
    .Y(_02676_)
  );
  NAND2X1 _09503_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_1_ ),
    .Y(_02677_)
  );
  NAND3X1 _09504_ (
    .A(execution_unit_0.register_file_0.r1_0_ ),
    .B(_02981_),
    .C(_02677_),
    .Y(_02678_)
  );
  NOR2X1 _09505_ (
    .A(_02674_),
    .B(_02678_),
    .Y(_02016_)
  );
  NOR2X1 _09506_ (
    .A(_03062_),
    .B(_02675_),
    .Y(_02679_)
  );
  OAI21X1 _09507_ (
    .A(execution_unit_0.register_file_0.r1_1_ ),
    .B(_02674_),
    .C(_02981_),
    .Y(_02680_)
  );
  AOI21X1 _09508_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_1_ ),
    .C(_02676_),
    .Y(_02681_)
  );
  OAI21X1 _09509_ (
    .A(_02679_),
    .B(_02680_),
    .C(_02681_),
    .Y(_02682_)
  );
  OAI21X1 _09510_ (
    .A(execution_unit_0.alu_0.alu_out_1_ ),
    .B(_02677_),
    .C(_02682_),
    .Y(_02683_)
  );
  INVX1 _09511_ (
    .A(_02683_),
    .Y(_02023_)
  );
  AOI21X1 _09512_ (
    .A(_03083_),
    .B(_02674_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02684_)
  );
  OAI21X1 _09513_ (
    .A(execution_unit_0.register_file_0.r1_2_ ),
    .B(_02674_),
    .C(_02684_),
    .Y(_02685_)
  );
  AOI21X1 _09514_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_2_ ),
    .C(_02676_),
    .Y(_02686_)
  );
  AOI22X1 _09515_ (
    .A(_02959_),
    .B(_02676_),
    .C(_02685_),
    .D(_02686_),
    .Y(_02024_)
  );
  AOI21X1 _09516_ (
    .A(_02961_),
    .B(_02675_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02687_)
  );
  OAI21X1 _09517_ (
    .A(_03104_),
    .B(_02675_),
    .C(_02687_),
    .Y(_02688_)
  );
  AOI21X1 _09518_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_3_ ),
    .C(_02676_),
    .Y(_02689_)
  );
  AOI22X1 _09519_ (
    .A(_02962_),
    .B(_02676_),
    .C(_02688_),
    .D(_02689_),
    .Y(_02025_)
  );
  AOI21X1 _09520_ (
    .A(_02964_),
    .B(_02675_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02690_)
  );
  OAI21X1 _09521_ (
    .A(_03122_),
    .B(_02675_),
    .C(_02690_),
    .Y(_02691_)
  );
  AOI21X1 _09522_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_4_ ),
    .C(_02676_),
    .Y(_02692_)
  );
  AOI22X1 _09523_ (
    .A(_02965_),
    .B(_02676_),
    .C(_02691_),
    .D(_02692_),
    .Y(_02026_)
  );
  NOR2X1 _09524_ (
    .A(_03140_),
    .B(_02675_),
    .Y(_02693_)
  );
  OAI21X1 _09525_ (
    .A(execution_unit_0.register_file_0.r1_5_ ),
    .B(_02674_),
    .C(_02981_),
    .Y(_02694_)
  );
  NAND2X1 _09526_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_5_ ),
    .Y(_02695_)
  );
  OAI21X1 _09527_ (
    .A(_02693_),
    .B(_02694_),
    .C(_02695_),
    .Y(_02696_)
  );
  NAND2X1 _09528_ (
    .A(_02677_),
    .B(_02696_),
    .Y(_02697_)
  );
  OAI21X1 _09529_ (
    .A(_02966_),
    .B(_02677_),
    .C(_02697_),
    .Y(_02027_)
  );
  AOI21X1 _09530_ (
    .A(_03157_),
    .B(_02674_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02698_)
  );
  OAI21X1 _09531_ (
    .A(execution_unit_0.register_file_0.r1_6_ ),
    .B(_02674_),
    .C(_02698_),
    .Y(_02699_)
  );
  AOI21X1 _09532_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_6_ ),
    .C(_02676_),
    .Y(_02700_)
  );
  AOI22X1 _09533_ (
    .A(_02967_),
    .B(_02676_),
    .C(_02699_),
    .D(_02700_),
    .Y(_02028_)
  );
  NOR2X1 _09534_ (
    .A(execution_unit_0.register_file_0.r1_7_ ),
    .B(_02674_),
    .Y(_02701_)
  );
  OAI21X1 _09535_ (
    .A(_03177_),
    .B(_02675_),
    .C(_02981_),
    .Y(_02702_)
  );
  NAND2X1 _09536_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_02703_)
  );
  OAI21X1 _09537_ (
    .A(_02701_),
    .B(_02702_),
    .C(_02703_),
    .Y(_02704_)
  );
  NAND2X1 _09538_ (
    .A(_02677_),
    .B(_02704_),
    .Y(_02705_)
  );
  OAI21X1 _09539_ (
    .A(_02968_),
    .B(_02677_),
    .C(_02705_),
    .Y(_02029_)
  );
  AOI21X1 _09540_ (
    .A(_02969_),
    .B(_02675_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02706_)
  );
  OAI21X1 _09541_ (
    .A(_03195_),
    .B(_02675_),
    .C(_02706_),
    .Y(_02707_)
  );
  AOI21X1 _09542_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_8_ ),
    .C(_02676_),
    .Y(_02708_)
  );
  AOI22X1 _09543_ (
    .A(_02982_),
    .B(_02676_),
    .C(_02707_),
    .D(_02708_),
    .Y(_02030_)
  );
  NOR2X1 _09544_ (
    .A(_03212_),
    .B(_02675_),
    .Y(_02709_)
  );
  OAI21X1 _09545_ (
    .A(execution_unit_0.register_file_0.r1_9_ ),
    .B(_02674_),
    .C(_02981_),
    .Y(_02710_)
  );
  NAND2X1 _09546_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_9_ ),
    .Y(_02711_)
  );
  OAI21X1 _09547_ (
    .A(_02709_),
    .B(_02710_),
    .C(_02711_),
    .Y(_02712_)
  );
  NAND2X1 _09548_ (
    .A(_02677_),
    .B(_02712_),
    .Y(_02713_)
  );
  OAI21X1 _09549_ (
    .A(_02983_),
    .B(_02677_),
    .C(_02713_),
    .Y(_02031_)
  );
  AOI21X1 _09550_ (
    .A(_03231_),
    .B(_02674_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02714_)
  );
  OAI21X1 _09551_ (
    .A(execution_unit_0.register_file_0.r1_10_ ),
    .B(_02674_),
    .C(_02714_),
    .Y(_02715_)
  );
  AOI21X1 _09552_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_10_ ),
    .C(_02676_),
    .Y(_02716_)
  );
  AOI22X1 _09553_ (
    .A(_02984_),
    .B(_02676_),
    .C(_02715_),
    .D(_02716_),
    .Y(_02017_)
  );
  AOI21X1 _09554_ (
    .A(_02970_),
    .B(_02675_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02717_)
  );
  OAI21X1 _09555_ (
    .A(_03249_),
    .B(_02675_),
    .C(_02717_),
    .Y(_02718_)
  );
  AOI21X1 _09556_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_11_ ),
    .C(_02676_),
    .Y(_02719_)
  );
  AOI22X1 _09557_ (
    .A(_02985_),
    .B(_02676_),
    .C(_02718_),
    .D(_02719_),
    .Y(_02018_)
  );
  NOR2X1 _09558_ (
    .A(_03267_),
    .B(_02675_),
    .Y(_02720_)
  );
  OAI21X1 _09559_ (
    .A(execution_unit_0.register_file_0.r1_12_ ),
    .B(_02674_),
    .C(_02981_),
    .Y(_02721_)
  );
  NAND2X1 _09560_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_12_ ),
    .Y(_02722_)
  );
  OAI21X1 _09561_ (
    .A(_02720_),
    .B(_02721_),
    .C(_02722_),
    .Y(_02723_)
  );
  NAND2X1 _09562_ (
    .A(_02677_),
    .B(_02723_),
    .Y(_02724_)
  );
  OAI21X1 _09563_ (
    .A(_02986_),
    .B(_02677_),
    .C(_02724_),
    .Y(_02019_)
  );
  AOI21X1 _09564_ (
    .A(_02971_),
    .B(_02675_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02725_)
  );
  OAI21X1 _09565_ (
    .A(_03285_),
    .B(_02675_),
    .C(_02725_),
    .Y(_02726_)
  );
  AOI21X1 _09566_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_13_ ),
    .C(_02676_),
    .Y(_02727_)
  );
  AOI22X1 _09567_ (
    .A(_02987_),
    .B(_02676_),
    .C(_02726_),
    .D(_02727_),
    .Y(_02020_)
  );
  AOI21X1 _09568_ (
    .A(_02973_),
    .B(_02675_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02728_)
  );
  OAI21X1 _09569_ (
    .A(_03303_),
    .B(_02675_),
    .C(_02728_),
    .Y(_02729_)
  );
  AOI21X1 _09570_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_14_ ),
    .C(_02676_),
    .Y(_02730_)
  );
  AOI22X1 _09571_ (
    .A(_02988_),
    .B(_02676_),
    .C(_02729_),
    .D(_02730_),
    .Y(_02021_)
  );
  AOI21X1 _09572_ (
    .A(_02975_),
    .B(_02675_),
    .C(execution_unit_0.reg_sp_wr ),
    .Y(_02731_)
  );
  OAI21X1 _09573_ (
    .A(_02165_),
    .B(_02675_),
    .C(_02731_),
    .Y(_02732_)
  );
  AOI21X1 _09574_ (
    .A(execution_unit_0.reg_sp_wr ),
    .B(dbg_0.UNUSED_eu_mab_15_ ),
    .C(_02676_),
    .Y(_02733_)
  );
  AOI22X1 _09575_ (
    .A(_02989_),
    .B(_02676_),
    .C(_02732_),
    .D(_02733_),
    .Y(_02022_)
  );
  AOI21X1 _09576_ (
    .A(execution_unit_0.reg_dest_wr ),
    .B(execution_unit_0.inst_dest_0_ ),
    .C(execution_unit_0.reg_pc_call ),
    .Y(_02734_)
  );
  INVX1 _09577_ (
    .A(_02734_),
    .Y(execution_unit_0.pc_sw_wr )
  );
  AOI22X1 _09578_ (
    .A(execution_unit_0.register_file_0.r9_0_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_0_ ),
    .Y(_02735_)
  );
  AOI22X1 _09579_ (
    .A(execution_unit_0.register_file_0.r12_0_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_0_ ),
    .Y(_02736_)
  );
  NAND2X1 _09580_ (
    .A(_02735_),
    .B(_02736_),
    .Y(_02737_)
  );
  AOI22X1 _09581_ (
    .A(execution_unit_0.register_file_0.r13_0_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_0_ ),
    .Y(_02738_)
  );
  AOI22X1 _09582_ (
    .A(execution_unit_0.register_file_0.r6_0_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_0_ ),
    .Y(_02739_)
  );
  NAND2X1 _09583_ (
    .A(_02738_),
    .B(_02739_),
    .Y(_02740_)
  );
  NOR2X1 _09584_ (
    .A(_02737_),
    .B(_02740_),
    .Y(_02741_)
  );
  AOI22X1 _09585_ (
    .A(execution_unit_0.register_file_0.r15_0_ ),
    .B(execution_unit_0.inst_dest_15_ ),
    .C(execution_unit_0.inst_dest_2_ ),
    .D(execution_unit_0.alu_0.status_0_ ),
    .Y(_02742_)
  );
  AOI22X1 _09586_ (
    .A(execution_unit_0.register_file_0.r11_0_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_0_ ),
    .Y(_02743_)
  );
  NAND2X1 _09587_ (
    .A(_02742_),
    .B(_02743_),
    .Y(_02744_)
  );
  AOI22X1 _09588_ (
    .A(execution_unit_0.register_file_0.r4_0_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_0_ ),
    .Y(_02745_)
  );
  AOI22X1 _09589_ (
    .A(execution_unit_0.register_file_0.r14_0_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_0_ ),
    .Y(_02746_)
  );
  NAND2X1 _09590_ (
    .A(_02745_),
    .B(_02746_),
    .Y(_02747_)
  );
  NOR2X1 _09591_ (
    .A(_02744_),
    .B(_02747_),
    .Y(_02748_)
  );
  NAND2X1 _09592_ (
    .A(_02741_),
    .B(_02748_),
    .Y(dbg_0.dbg_reg_din_0_ )
  );
  AOI22X1 _09593_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_1_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_1_ ),
    .Y(_02749_)
  );
  AOI22X1 _09594_ (
    .A(execution_unit_0.register_file_0.r3_1_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_1_ ),
    .Y(_02750_)
  );
  NAND2X1 _09595_ (
    .A(_02749_),
    .B(_02750_),
    .Y(_02751_)
  );
  AOI22X1 _09596_ (
    .A(execution_unit_0.register_file_0.r6_1_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_2_ ),
    .D(execution_unit_0.alu_0.status_1_ ),
    .Y(_02752_)
  );
  AOI22X1 _09597_ (
    .A(execution_unit_0.register_file_0.r10_1_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_1_ ),
    .Y(_02753_)
  );
  NAND2X1 _09598_ (
    .A(_02752_),
    .B(_02753_),
    .Y(_02754_)
  );
  NOR2X1 _09599_ (
    .A(_02751_),
    .B(_02754_),
    .Y(_02755_)
  );
  AOI22X1 _09600_ (
    .A(execution_unit_0.register_file_0.r14_1_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_1_ ),
    .Y(_02756_)
  );
  AOI22X1 _09601_ (
    .A(execution_unit_0.register_file_0.r13_1_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_1_ ),
    .Y(_02757_)
  );
  NAND2X1 _09602_ (
    .A(_02756_),
    .B(_02757_),
    .Y(_02758_)
  );
  AOI22X1 _09603_ (
    .A(execution_unit_0.register_file_0.r12_1_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_1_ ),
    .Y(_02759_)
  );
  AOI22X1 _09604_ (
    .A(execution_unit_0.register_file_0.r9_1_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_1_ ),
    .Y(_02760_)
  );
  NAND2X1 _09605_ (
    .A(_02759_),
    .B(_02760_),
    .Y(_02761_)
  );
  NOR2X1 _09606_ (
    .A(_02758_),
    .B(_02761_),
    .Y(_02762_)
  );
  NAND2X1 _09607_ (
    .A(_02755_),
    .B(_02762_),
    .Y(dbg_0.dbg_reg_din_1_ )
  );
  AOI22X1 _09608_ (
    .A(execution_unit_0.register_file_0.r14_2_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_2_ ),
    .Y(_02763_)
  );
  AOI22X1 _09609_ (
    .A(execution_unit_0.register_file_0.r10_2_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_2_ ),
    .Y(_02764_)
  );
  NAND2X1 _09610_ (
    .A(_02763_),
    .B(_02764_),
    .Y(_02765_)
  );
  AOI22X1 _09611_ (
    .A(execution_unit_0.register_file_0.r1_2_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_2_ ),
    .Y(_02766_)
  );
  AOI22X1 _09612_ (
    .A(execution_unit_0.register_file_0.r13_2_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_2_ ),
    .Y(_02767_)
  );
  NAND2X1 _09613_ (
    .A(_02766_),
    .B(_02767_),
    .Y(_02768_)
  );
  NOR2X1 _09614_ (
    .A(_02765_),
    .B(_02768_),
    .Y(_02769_)
  );
  AOI22X1 _09615_ (
    .A(execution_unit_0.register_file_0.r5_2_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_2_ ),
    .D(execution_unit_0.alu_0.status_2_ ),
    .Y(_02770_)
  );
  AOI22X1 _09616_ (
    .A(execution_unit_0.register_file_0.r9_2_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_2_ ),
    .Y(_02771_)
  );
  AOI22X1 _09617_ (
    .A(execution_unit_0.register_file_0.r6_2_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_2_ ),
    .Y(_02772_)
  );
  NAND2X1 _09618_ (
    .A(_02771_),
    .B(_02772_),
    .Y(_02773_)
  );
  AOI22X1 _09619_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_2_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_2_ ),
    .Y(_02774_)
  );
  NAND2X1 _09620_ (
    .A(_02770_),
    .B(_02774_),
    .Y(_02775_)
  );
  NOR2X1 _09621_ (
    .A(_02773_),
    .B(_02775_),
    .Y(_02776_)
  );
  NAND2X1 _09622_ (
    .A(_02769_),
    .B(_02776_),
    .Y(dbg_0.dbg_reg_din_2_ )
  );
  AOI22X1 _09623_ (
    .A(execution_unit_0.register_file_0.r4_3_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_3_ ),
    .Y(_02777_)
  );
  AOI22X1 _09624_ (
    .A(execution_unit_0.register_file_0.r14_3_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_3_ ),
    .Y(_02778_)
  );
  NAND2X1 _09625_ (
    .A(_02777_),
    .B(_02778_),
    .Y(_02779_)
  );
  AOI22X1 _09626_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_3_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_3_ ),
    .Y(_02780_)
  );
  AOI22X1 _09627_ (
    .A(execution_unit_0.register_file_0.r6_3_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_3_ ),
    .Y(_02781_)
  );
  NAND2X1 _09628_ (
    .A(_02780_),
    .B(_02781_),
    .Y(_02782_)
  );
  NOR2X1 _09629_ (
    .A(_02779_),
    .B(_02782_),
    .Y(_02783_)
  );
  AOI22X1 _09630_ (
    .A(execution_unit_0.register_file_0.r13_3_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_3_ ),
    .Y(_02784_)
  );
  AOI22X1 _09631_ (
    .A(execution_unit_0.register_file_0.r11_3_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_3_ ),
    .Y(_02785_)
  );
  NAND2X1 _09632_ (
    .A(_02784_),
    .B(_02785_),
    .Y(_02786_)
  );
  AOI22X1 _09633_ (
    .A(execution_unit_0.register_file_0.r10_3_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_2_ ),
    .D(execution_unit_0.gie ),
    .Y(_02787_)
  );
  AOI22X1 _09634_ (
    .A(execution_unit_0.register_file_0.r12_3_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_3_ ),
    .Y(_02788_)
  );
  NAND2X1 _09635_ (
    .A(_02787_),
    .B(_02788_),
    .Y(_02789_)
  );
  NOR2X1 _09636_ (
    .A(_02786_),
    .B(_02789_),
    .Y(_02790_)
  );
  NAND2X1 _09637_ (
    .A(_02783_),
    .B(_02790_),
    .Y(dbg_0.dbg_reg_din_3_ )
  );
  AOI22X1 _09638_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_4_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_4_ ),
    .Y(_02791_)
  );
  AOI22X1 _09639_ (
    .A(execution_unit_0.register_file_0.r9_4_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_4_ ),
    .Y(_02792_)
  );
  NAND2X1 _09640_ (
    .A(_02791_),
    .B(_02792_),
    .Y(_02793_)
  );
  AOI22X1 _09641_ (
    .A(execution_unit_0.register_file_0.r13_4_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_4_ ),
    .Y(_02794_)
  );
  AOI22X1 _09642_ (
    .A(execution_unit_0.register_file_0.r12_4_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_4_ ),
    .Y(_02795_)
  );
  NAND2X1 _09643_ (
    .A(_02794_),
    .B(_02795_),
    .Y(_02796_)
  );
  NOR2X1 _09644_ (
    .A(_02793_),
    .B(_02796_),
    .Y(_02797_)
  );
  AOI22X1 _09645_ (
    .A(execution_unit_0.register_file_0.r10_4_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_4_ ),
    .Y(_02798_)
  );
  AOI22X1 _09646_ (
    .A(execution_unit_0.register_file_0.r3_4_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_2_ ),
    .D(execution_unit_0.register_file_0.r2_4_ ),
    .Y(_02799_)
  );
  NAND2X1 _09647_ (
    .A(_02798_),
    .B(_02799_),
    .Y(_02800_)
  );
  AOI22X1 _09648_ (
    .A(execution_unit_0.register_file_0.r14_4_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_4_ ),
    .Y(_02801_)
  );
  AOI22X1 _09649_ (
    .A(execution_unit_0.register_file_0.r8_4_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_4_ ),
    .Y(_02802_)
  );
  NAND2X1 _09650_ (
    .A(_02801_),
    .B(_02802_),
    .Y(_02803_)
  );
  NOR2X1 _09651_ (
    .A(_02800_),
    .B(_02803_),
    .Y(_02804_)
  );
  NAND2X1 _09652_ (
    .A(_02797_),
    .B(_02804_),
    .Y(dbg_0.dbg_reg_din_4_ )
  );
  AOI22X1 _09653_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_5_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_5_ ),
    .Y(_02805_)
  );
  AOI22X1 _09654_ (
    .A(execution_unit_0.register_file_0.r6_5_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_2_ ),
    .D(clock_module_0.oscoff ),
    .Y(_02806_)
  );
  NAND2X1 _09655_ (
    .A(_02805_),
    .B(_02806_),
    .Y(_02807_)
  );
  AOI22X1 _09656_ (
    .A(execution_unit_0.register_file_0.r3_5_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_5_ ),
    .Y(_02808_)
  );
  AOI22X1 _09657_ (
    .A(execution_unit_0.register_file_0.r8_5_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_5_ ),
    .Y(_02809_)
  );
  NAND2X1 _09658_ (
    .A(_02808_),
    .B(_02809_),
    .Y(_02810_)
  );
  NOR2X1 _09659_ (
    .A(_02807_),
    .B(_02810_),
    .Y(_02811_)
  );
  AOI22X1 _09660_ (
    .A(execution_unit_0.register_file_0.r11_5_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_5_ ),
    .Y(_02812_)
  );
  AOI22X1 _09661_ (
    .A(execution_unit_0.register_file_0.r14_5_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_5_ ),
    .Y(_02813_)
  );
  NAND2X1 _09662_ (
    .A(_02812_),
    .B(_02813_),
    .Y(_02814_)
  );
  AOI22X1 _09663_ (
    .A(execution_unit_0.register_file_0.r13_5_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_5_ ),
    .Y(_02815_)
  );
  AOI22X1 _09664_ (
    .A(execution_unit_0.register_file_0.r5_5_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_5_ ),
    .Y(_02816_)
  );
  NAND2X1 _09665_ (
    .A(_02815_),
    .B(_02816_),
    .Y(_02817_)
  );
  NOR2X1 _09666_ (
    .A(_02814_),
    .B(_02817_),
    .Y(_02818_)
  );
  NAND2X1 _09667_ (
    .A(_02811_),
    .B(_02818_),
    .Y(dbg_0.dbg_reg_din_5_ )
  );
  NAND2X1 _09668_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_6_ ),
    .Y(_02819_)
  );
  NAND2X1 _09669_ (
    .A(execution_unit_0.register_file_0.r4_6_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .Y(_02820_)
  );
  AOI22X1 _09670_ (
    .A(execution_unit_0.register_file_0.r7_6_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_6_ ),
    .Y(_02821_)
  );
  AOI22X1 _09671_ (
    .A(execution_unit_0.register_file_0.r10_6_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_6_ ),
    .Y(_02822_)
  );
  AOI22X1 _09672_ (
    .A(execution_unit_0.register_file_0.r12_6_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_6_ ),
    .Y(_02823_)
  );
  NAND2X1 _09673_ (
    .A(_02822_),
    .B(_02823_),
    .Y(_02824_)
  );
  AOI21X1 _09674_ (
    .A(execution_unit_0.register_file_0.r14_6_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(_02824_),
    .Y(_02825_)
  );
  NAND3X1 _09675_ (
    .A(_02819_),
    .B(_02820_),
    .C(_02821_),
    .Y(_02826_)
  );
  AOI22X1 _09676_ (
    .A(execution_unit_0.register_file_0.r9_6_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_6_ ),
    .Y(_02827_)
  );
  AOI22X1 _09677_ (
    .A(execution_unit_0.register_file_0.r11_6_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_6_ ),
    .Y(_02828_)
  );
  AOI22X1 _09678_ (
    .A(execution_unit_0.register_file_0.r13_6_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_6_ ),
    .Y(_02829_)
  );
  NAND3X1 _09679_ (
    .A(_02827_),
    .B(_02828_),
    .C(_02829_),
    .Y(_02830_)
  );
  NOR2X1 _09680_ (
    .A(_02826_),
    .B(_02830_),
    .Y(_02831_)
  );
  NAND2X1 _09681_ (
    .A(_02825_),
    .B(_02831_),
    .Y(dbg_0.dbg_reg_din_6_ )
  );
  AOI22X1 _09682_ (
    .A(execution_unit_0.register_file_0.r8_7_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_7_ ),
    .Y(_02832_)
  );
  AOI22X1 _09683_ (
    .A(execution_unit_0.register_file_0.r10_7_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_7_ ),
    .Y(_02833_)
  );
  NAND2X1 _09684_ (
    .A(_02832_),
    .B(_02833_),
    .Y(_02834_)
  );
  AOI22X1 _09685_ (
    .A(execution_unit_0.register_file_0.r11_7_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_7_ ),
    .Y(_02835_)
  );
  AOI22X1 _09686_ (
    .A(execution_unit_0.register_file_0.r14_7_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_7_ ),
    .Y(_02836_)
  );
  NAND2X1 _09687_ (
    .A(_02835_),
    .B(_02836_),
    .Y(_02837_)
  );
  NOR2X1 _09688_ (
    .A(_02834_),
    .B(_02837_),
    .Y(_02838_)
  );
  AOI22X1 _09689_ (
    .A(execution_unit_0.register_file_0.r13_7_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_2_ ),
    .D(clock_module_0.scg1 ),
    .Y(_02839_)
  );
  AOI22X1 _09690_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_7_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_7_ ),
    .Y(_02840_)
  );
  NAND2X1 _09691_ (
    .A(_02839_),
    .B(_02840_),
    .Y(_02841_)
  );
  AOI22X1 _09692_ (
    .A(execution_unit_0.register_file_0.r4_7_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_7_ ),
    .Y(_02842_)
  );
  AOI22X1 _09693_ (
    .A(execution_unit_0.register_file_0.r9_7_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_7_ ),
    .Y(_02843_)
  );
  NAND2X1 _09694_ (
    .A(_02842_),
    .B(_02843_),
    .Y(_02844_)
  );
  NOR2X1 _09695_ (
    .A(_02841_),
    .B(_02844_),
    .Y(_02845_)
  );
  NAND2X1 _09696_ (
    .A(_02838_),
    .B(_02845_),
    .Y(dbg_0.dbg_reg_din_7_ )
  );
  AOI22X1 _09697_ (
    .A(execution_unit_0.register_file_0.r8_8_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_8_ ),
    .Y(_02846_)
  );
  AOI22X1 _09698_ (
    .A(execution_unit_0.register_file_0.r10_8_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_8_ ),
    .Y(_02847_)
  );
  NAND2X1 _09699_ (
    .A(_02846_),
    .B(_02847_),
    .Y(_02848_)
  );
  AOI22X1 _09700_ (
    .A(execution_unit_0.register_file_0.r12_8_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_8_ ),
    .Y(_02849_)
  );
  AOI22X1 _09701_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_8_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_8_ ),
    .Y(_02850_)
  );
  NAND2X1 _09702_ (
    .A(_02849_),
    .B(_02850_),
    .Y(_02851_)
  );
  NOR2X1 _09703_ (
    .A(_02848_),
    .B(_02851_),
    .Y(_02852_)
  );
  AOI22X1 _09704_ (
    .A(execution_unit_0.register_file_0.r6_8_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_8_ ),
    .Y(_02853_)
  );
  AOI22X1 _09705_ (
    .A(execution_unit_0.register_file_0.r7_8_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_2_ ),
    .D(execution_unit_0.alu_0.status_3_ ),
    .Y(_02854_)
  );
  NAND2X1 _09706_ (
    .A(_02853_),
    .B(_02854_),
    .Y(_02855_)
  );
  AOI22X1 _09707_ (
    .A(execution_unit_0.register_file_0.r14_8_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_8_ ),
    .Y(_02856_)
  );
  AOI22X1 _09708_ (
    .A(execution_unit_0.register_file_0.r13_8_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_8_ ),
    .Y(_02857_)
  );
  NAND2X1 _09709_ (
    .A(_02856_),
    .B(_02857_),
    .Y(_02858_)
  );
  NOR2X1 _09710_ (
    .A(_02855_),
    .B(_02858_),
    .Y(_02859_)
  );
  NAND2X1 _09711_ (
    .A(_02852_),
    .B(_02859_),
    .Y(dbg_0.dbg_reg_din_8_ )
  );
  NAND2X1 _09712_ (
    .A(execution_unit_0.register_file_0.r1_9_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .Y(_02860_)
  );
  NAND2X1 _09713_ (
    .A(execution_unit_0.register_file_0.r5_9_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .Y(_02861_)
  );
  AOI22X1 _09714_ (
    .A(execution_unit_0.register_file_0.r14_9_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_9_ ),
    .Y(_02862_)
  );
  AOI22X1 _09715_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_9_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_9_ ),
    .Y(_02863_)
  );
  NAND2X1 _09716_ (
    .A(_02862_),
    .B(_02863_),
    .Y(_02864_)
  );
  AOI21X1 _09717_ (
    .A(execution_unit_0.register_file_0.r3_9_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(_02864_),
    .Y(_02865_)
  );
  AOI22X1 _09718_ (
    .A(execution_unit_0.register_file_0.r10_9_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_9_ ),
    .Y(_02866_)
  );
  NAND3X1 _09719_ (
    .A(_02860_),
    .B(_02861_),
    .C(_02866_),
    .Y(_02867_)
  );
  AOI22X1 _09720_ (
    .A(execution_unit_0.register_file_0.r7_9_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_9_ ),
    .Y(_02868_)
  );
  AOI22X1 _09721_ (
    .A(execution_unit_0.register_file_0.r11_9_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_9_ ),
    .Y(_02869_)
  );
  AOI22X1 _09722_ (
    .A(execution_unit_0.register_file_0.r13_9_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_9_ ),
    .Y(_02870_)
  );
  NAND3X1 _09723_ (
    .A(_02868_),
    .B(_02869_),
    .C(_02870_),
    .Y(_02871_)
  );
  NOR2X1 _09724_ (
    .A(_02867_),
    .B(_02871_),
    .Y(_02872_)
  );
  NAND2X1 _09725_ (
    .A(_02865_),
    .B(_02872_),
    .Y(dbg_0.dbg_reg_din_9_ )
  );
  AOI22X1 _09726_ (
    .A(execution_unit_0.register_file_0.r10_10_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_10_ ),
    .Y(_02873_)
  );
  NAND2X1 _09727_ (
    .A(execution_unit_0.register_file_0.r1_10_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .Y(_02874_)
  );
  NAND2X1 _09728_ (
    .A(execution_unit_0.register_file_0.r5_10_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .Y(_02875_)
  );
  AOI22X1 _09729_ (
    .A(execution_unit_0.register_file_0.r9_10_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_8_ ),
    .D(execution_unit_0.register_file_0.r8_10_ ),
    .Y(_02876_)
  );
  NAND2X1 _09730_ (
    .A(_02875_),
    .B(_02876_),
    .Y(_02877_)
  );
  AOI21X1 _09731_ (
    .A(dbg_0.UNUSED_pc_10_ ),
    .B(execution_unit_0.inst_dest_0_ ),
    .C(_02877_),
    .Y(_02878_)
  );
  AOI22X1 _09732_ (
    .A(execution_unit_0.register_file_0.r14_10_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_10_ ),
    .Y(_02879_)
  );
  NAND2X1 _09733_ (
    .A(_02873_),
    .B(_02879_),
    .Y(_02880_)
  );
  AOI21X1 _09734_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_10_ ),
    .C(_02880_),
    .Y(_02881_)
  );
  AOI22X1 _09735_ (
    .A(execution_unit_0.register_file_0.r11_10_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_10_ ),
    .Y(_02882_)
  );
  AOI22X1 _09736_ (
    .A(execution_unit_0.register_file_0.r13_10_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_10_ ),
    .Y(_02883_)
  );
  NAND3X1 _09737_ (
    .A(_02874_),
    .B(_02882_),
    .C(_02883_),
    .Y(_02884_)
  );
  AOI21X1 _09738_ (
    .A(execution_unit_0.register_file_0.r7_10_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(_02884_),
    .Y(_02885_)
  );
  NAND3X1 _09739_ (
    .A(_02878_),
    .B(_02881_),
    .C(_02885_),
    .Y(dbg_0.dbg_reg_din_10_ )
  );
  NAND2X1 _09740_ (
    .A(execution_unit_0.register_file_0.r13_11_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .Y(_02886_)
  );
  NAND2X1 _09741_ (
    .A(dbg_0.UNUSED_pc_11_ ),
    .B(execution_unit_0.inst_dest_0_ ),
    .Y(_02887_)
  );
  AOI22X1 _09742_ (
    .A(execution_unit_0.register_file_0.r12_11_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_11_ ),
    .Y(_02888_)
  );
  AOI22X1 _09743_ (
    .A(execution_unit_0.register_file_0.r10_11_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_11_ ),
    .Y(_02889_)
  );
  NAND2X1 _09744_ (
    .A(_02887_),
    .B(_02889_),
    .Y(_02890_)
  );
  AOI22X1 _09745_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_11_ ),
    .C(execution_unit_0.inst_dest_14_ ),
    .D(execution_unit_0.register_file_0.r14_11_ ),
    .Y(_02891_)
  );
  NAND2X1 _09746_ (
    .A(_02886_),
    .B(_02891_),
    .Y(_02892_)
  );
  NOR2X1 _09747_ (
    .A(_02890_),
    .B(_02892_),
    .Y(_02893_)
  );
  AOI22X1 _09748_ (
    .A(execution_unit_0.register_file_0.r11_11_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_11_ ),
    .Y(_02894_)
  );
  AOI22X1 _09749_ (
    .A(execution_unit_0.register_file_0.r9_11_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_11_ ),
    .Y(_02895_)
  );
  AOI22X1 _09750_ (
    .A(execution_unit_0.register_file_0.r8_11_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_11_ ),
    .Y(_02896_)
  );
  NAND3X1 _09751_ (
    .A(_02894_),
    .B(_02895_),
    .C(_02896_),
    .Y(_02897_)
  );
  AOI21X1 _09752_ (
    .A(execution_unit_0.register_file_0.r3_11_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(_02897_),
    .Y(_02898_)
  );
  NAND3X1 _09753_ (
    .A(_02888_),
    .B(_02893_),
    .C(_02898_),
    .Y(dbg_0.dbg_reg_din_11_ )
  );
  NAND2X1 _09754_ (
    .A(execution_unit_0.register_file_0.r1_12_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .Y(_02899_)
  );
  AOI22X1 _09755_ (
    .A(execution_unit_0.register_file_0.r11_12_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_12_ ),
    .Y(_02900_)
  );
  NAND2X1 _09756_ (
    .A(execution_unit_0.register_file_0.r5_12_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .Y(_02901_)
  );
  AOI22X1 _09757_ (
    .A(execution_unit_0.register_file_0.r13_12_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_12_ ),
    .Y(_02902_)
  );
  AOI22X1 _09758_ (
    .A(execution_unit_0.register_file_0.r14_12_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_12_ ),
    .D(execution_unit_0.register_file_0.r12_12_ ),
    .Y(_02903_)
  );
  AOI22X1 _09759_ (
    .A(execution_unit_0.register_file_0.r10_12_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_12_ ),
    .Y(_02904_)
  );
  NAND2X1 _09760_ (
    .A(_02903_),
    .B(_02904_),
    .Y(_02905_)
  );
  AOI21X1 _09761_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_12_ ),
    .C(_02905_),
    .Y(_02906_)
  );
  AOI22X1 _09762_ (
    .A(execution_unit_0.register_file_0.r8_12_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_7_ ),
    .D(execution_unit_0.register_file_0.r7_12_ ),
    .Y(_02907_)
  );
  NAND3X1 _09763_ (
    .A(_02899_),
    .B(_02901_),
    .C(_02907_),
    .Y(_02908_)
  );
  AOI22X1 _09764_ (
    .A(execution_unit_0.register_file_0.r9_12_ ),
    .B(execution_unit_0.inst_dest_9_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_12_ ),
    .Y(_02909_)
  );
  NAND3X1 _09765_ (
    .A(_02900_),
    .B(_02902_),
    .C(_02909_),
    .Y(_02910_)
  );
  NOR2X1 _09766_ (
    .A(_02908_),
    .B(_02910_),
    .Y(_02911_)
  );
  NAND2X1 _09767_ (
    .A(_02906_),
    .B(_02911_),
    .Y(dbg_0.dbg_reg_din_12_ )
  );
  AOI22X1 _09768_ (
    .A(execution_unit_0.register_file_0.r7_13_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_13_ ),
    .Y(_02912_)
  );
  AOI22X1 _09769_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_13_ ),
    .C(execution_unit_0.inst_dest_13_ ),
    .D(execution_unit_0.register_file_0.r13_13_ ),
    .Y(_02913_)
  );
  AOI22X1 _09770_ (
    .A(execution_unit_0.register_file_0.r14_13_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_13_ ),
    .Y(_02914_)
  );
  AOI22X1 _09771_ (
    .A(execution_unit_0.register_file_0.r8_13_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_13_ ),
    .Y(_02915_)
  );
  AND2X1 _09772_ (
    .A(_02914_),
    .B(_02915_),
    .Y(_02916_)
  );
  NAND3X1 _09773_ (
    .A(_02912_),
    .B(_02913_),
    .C(_02916_),
    .Y(_02917_)
  );
  AOI22X1 _09774_ (
    .A(execution_unit_0.register_file_0.r4_13_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_13_ ),
    .Y(_02918_)
  );
  INVX1 _09775_ (
    .A(_02918_),
    .Y(_02919_)
  );
  AOI21X1 _09776_ (
    .A(execution_unit_0.register_file_0.r10_13_ ),
    .B(execution_unit_0.inst_dest_10_ ),
    .C(_02919_),
    .Y(_02920_)
  );
  AOI22X1 _09777_ (
    .A(execution_unit_0.register_file_0.r11_13_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .C(execution_unit_0.inst_dest_6_ ),
    .D(execution_unit_0.register_file_0.r6_13_ ),
    .Y(_02921_)
  );
  AOI22X1 _09778_ (
    .A(execution_unit_0.register_file_0.r12_13_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_13_ ),
    .Y(_02922_)
  );
  NAND3X1 _09779_ (
    .A(_02920_),
    .B(_02921_),
    .C(_02922_),
    .Y(_02923_)
  );
  OR2X1 _09780_ (
    .A(_02917_),
    .B(_02923_),
    .Y(dbg_0.dbg_reg_din_13_ )
  );
  NAND2X1 _09781_ (
    .A(execution_unit_0.register_file_0.r7_14_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .Y(_02924_)
  );
  AOI22X1 _09782_ (
    .A(execution_unit_0.register_file_0.r6_14_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_1_ ),
    .D(execution_unit_0.register_file_0.r1_14_ ),
    .Y(_02925_)
  );
  AOI22X1 _09783_ (
    .A(execution_unit_0.register_file_0.r5_14_ ),
    .B(execution_unit_0.inst_dest_5_ ),
    .C(execution_unit_0.inst_dest_3_ ),
    .D(execution_unit_0.register_file_0.r3_14_ ),
    .Y(_02926_)
  );
  AOI22X1 _09784_ (
    .A(execution_unit_0.register_file_0.r8_14_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(execution_unit_0.inst_dest_4_ ),
    .D(execution_unit_0.register_file_0.r4_14_ ),
    .Y(_02927_)
  );
  OAI21X1 _09785_ (
    .A(_02972_),
    .B(_02976_),
    .C(_02927_),
    .Y(_02928_)
  );
  AOI21X1 _09786_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_14_ ),
    .C(_02928_),
    .Y(_02929_)
  );
  AOI22X1 _09787_ (
    .A(execution_unit_0.register_file_0.r12_14_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_11_ ),
    .D(execution_unit_0.register_file_0.r11_14_ ),
    .Y(_02930_)
  );
  AOI22X1 _09788_ (
    .A(execution_unit_0.register_file_0.r13_14_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_14_ ),
    .Y(_02931_)
  );
  NAND2X1 _09789_ (
    .A(_02930_),
    .B(_02931_),
    .Y(_02932_)
  );
  AOI21X1 _09790_ (
    .A(execution_unit_0.register_file_0.r14_14_ ),
    .B(execution_unit_0.inst_dest_14_ ),
    .C(_02932_),
    .Y(_02933_)
  );
  NAND3X1 _09791_ (
    .A(_02924_),
    .B(_02925_),
    .C(_02926_),
    .Y(_02934_)
  );
  AOI21X1 _09792_ (
    .A(dbg_0.UNUSED_pc_14_ ),
    .B(execution_unit_0.inst_dest_0_ ),
    .C(_02934_),
    .Y(_02935_)
  );
  NAND3X1 _09793_ (
    .A(_02929_),
    .B(_02933_),
    .C(_02935_),
    .Y(dbg_0.dbg_reg_din_14_ )
  );
  NAND2X1 _09794_ (
    .A(execution_unit_0.register_file_0.r11_15_ ),
    .B(execution_unit_0.inst_dest_11_ ),
    .Y(_02936_)
  );
  NAND2X1 _09795_ (
    .A(execution_unit_0.register_file_0.r4_15_ ),
    .B(execution_unit_0.inst_dest_4_ ),
    .Y(_02937_)
  );
  AOI22X1 _09796_ (
    .A(execution_unit_0.inst_dest_15_ ),
    .B(execution_unit_0.register_file_0.r15_15_ ),
    .C(execution_unit_0.register_file_0.r14_15_ ),
    .D(execution_unit_0.inst_dest_14_ ),
    .Y(_02938_)
  );
  NAND2X1 _09797_ (
    .A(_02937_),
    .B(_02938_),
    .Y(_02939_)
  );
  AOI21X1 _09798_ (
    .A(execution_unit_0.register_file_0.r7_15_ ),
    .B(execution_unit_0.inst_dest_7_ ),
    .C(_02939_),
    .Y(_02940_)
  );
  AOI22X1 _09799_ (
    .A(execution_unit_0.register_file_0.r1_15_ ),
    .B(execution_unit_0.inst_dest_1_ ),
    .C(execution_unit_0.inst_dest_0_ ),
    .D(dbg_0.UNUSED_pc_15_ ),
    .Y(_02941_)
  );
  AOI22X1 _09800_ (
    .A(execution_unit_0.register_file_0.r6_15_ ),
    .B(execution_unit_0.inst_dest_6_ ),
    .C(execution_unit_0.inst_dest_5_ ),
    .D(execution_unit_0.register_file_0.r5_15_ ),
    .Y(_02942_)
  );
  NAND2X1 _09801_ (
    .A(_02941_),
    .B(_02942_),
    .Y(_02943_)
  );
  AOI21X1 _09802_ (
    .A(execution_unit_0.register_file_0.r3_15_ ),
    .B(execution_unit_0.inst_dest_3_ ),
    .C(_02943_),
    .Y(_02944_)
  );
  AOI22X1 _09803_ (
    .A(execution_unit_0.register_file_0.r13_15_ ),
    .B(execution_unit_0.inst_dest_13_ ),
    .C(execution_unit_0.inst_dest_10_ ),
    .D(execution_unit_0.register_file_0.r10_15_ ),
    .Y(_02945_)
  );
  AOI22X1 _09804_ (
    .A(execution_unit_0.register_file_0.r12_15_ ),
    .B(execution_unit_0.inst_dest_12_ ),
    .C(execution_unit_0.inst_dest_9_ ),
    .D(execution_unit_0.register_file_0.r9_15_ ),
    .Y(_02946_)
  );
  NAND3X1 _09805_ (
    .A(_02936_),
    .B(_02945_),
    .C(_02946_),
    .Y(_02947_)
  );
  AOI21X1 _09806_ (
    .A(execution_unit_0.register_file_0.r8_15_ ),
    .B(execution_unit_0.inst_dest_8_ ),
    .C(_02947_),
    .Y(_02948_)
  );
  NAND3X1 _09807_ (
    .A(_02940_),
    .B(_02944_),
    .C(_02948_),
    .Y(dbg_0.dbg_reg_din_15_ )
  );
  DFFSR _09808_ (
    .CLK(dco_clk),
    .D(_02000_),
    .Q(execution_unit_0.register_file_0.r15_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09809_ (
    .CLK(dco_clk),
    .D(_02007_),
    .Q(execution_unit_0.register_file_0.r15_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09810_ (
    .CLK(dco_clk),
    .D(_02008_),
    .Q(execution_unit_0.register_file_0.r15_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09811_ (
    .CLK(dco_clk),
    .D(_02009_),
    .Q(execution_unit_0.register_file_0.r15_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09812_ (
    .CLK(dco_clk),
    .D(_02010_),
    .Q(execution_unit_0.register_file_0.r15_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09813_ (
    .CLK(dco_clk),
    .D(_02011_),
    .Q(execution_unit_0.register_file_0.r15_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09814_ (
    .CLK(dco_clk),
    .D(_02012_),
    .Q(execution_unit_0.register_file_0.r15_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09815_ (
    .CLK(dco_clk),
    .D(_02013_),
    .Q(execution_unit_0.register_file_0.r15_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09816_ (
    .CLK(dco_clk),
    .D(_02014_),
    .Q(execution_unit_0.register_file_0.r15_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09817_ (
    .CLK(dco_clk),
    .D(_02015_),
    .Q(execution_unit_0.register_file_0.r15_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09818_ (
    .CLK(dco_clk),
    .D(_02001_),
    .Q(execution_unit_0.register_file_0.r15_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09819_ (
    .CLK(dco_clk),
    .D(_02002_),
    .Q(execution_unit_0.register_file_0.r15_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09820_ (
    .CLK(dco_clk),
    .D(_02003_),
    .Q(execution_unit_0.register_file_0.r15_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09821_ (
    .CLK(dco_clk),
    .D(_02004_),
    .Q(execution_unit_0.register_file_0.r15_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09822_ (
    .CLK(dco_clk),
    .D(_02005_),
    .Q(execution_unit_0.register_file_0.r15_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09823_ (
    .CLK(dco_clk),
    .D(_02006_),
    .Q(execution_unit_0.register_file_0.r15_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09824_ (
    .CLK(dco_clk),
    .D(_01984_),
    .Q(execution_unit_0.register_file_0.r14_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09825_ (
    .CLK(dco_clk),
    .D(_01991_),
    .Q(execution_unit_0.register_file_0.r14_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09826_ (
    .CLK(dco_clk),
    .D(_01992_),
    .Q(execution_unit_0.register_file_0.r14_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09827_ (
    .CLK(dco_clk),
    .D(_01993_),
    .Q(execution_unit_0.register_file_0.r14_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09828_ (
    .CLK(dco_clk),
    .D(_01994_),
    .Q(execution_unit_0.register_file_0.r14_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09829_ (
    .CLK(dco_clk),
    .D(_01995_),
    .Q(execution_unit_0.register_file_0.r14_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09830_ (
    .CLK(dco_clk),
    .D(_01996_),
    .Q(execution_unit_0.register_file_0.r14_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09831_ (
    .CLK(dco_clk),
    .D(_01997_),
    .Q(execution_unit_0.register_file_0.r14_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09832_ (
    .CLK(dco_clk),
    .D(_01998_),
    .Q(execution_unit_0.register_file_0.r14_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09833_ (
    .CLK(dco_clk),
    .D(_01999_),
    .Q(execution_unit_0.register_file_0.r14_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09834_ (
    .CLK(dco_clk),
    .D(_01985_),
    .Q(execution_unit_0.register_file_0.r14_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09835_ (
    .CLK(dco_clk),
    .D(_01986_),
    .Q(execution_unit_0.register_file_0.r14_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09836_ (
    .CLK(dco_clk),
    .D(_01987_),
    .Q(execution_unit_0.register_file_0.r14_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09837_ (
    .CLK(dco_clk),
    .D(_01988_),
    .Q(execution_unit_0.register_file_0.r14_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09838_ (
    .CLK(dco_clk),
    .D(_01989_),
    .Q(execution_unit_0.register_file_0.r14_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09839_ (
    .CLK(dco_clk),
    .D(_01990_),
    .Q(execution_unit_0.register_file_0.r14_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09840_ (
    .CLK(dco_clk),
    .D(_01968_),
    .Q(execution_unit_0.register_file_0.r13_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09841_ (
    .CLK(dco_clk),
    .D(_01975_),
    .Q(execution_unit_0.register_file_0.r13_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09842_ (
    .CLK(dco_clk),
    .D(_01976_),
    .Q(execution_unit_0.register_file_0.r13_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09843_ (
    .CLK(dco_clk),
    .D(_01977_),
    .Q(execution_unit_0.register_file_0.r13_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09844_ (
    .CLK(dco_clk),
    .D(_01978_),
    .Q(execution_unit_0.register_file_0.r13_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09845_ (
    .CLK(dco_clk),
    .D(_01979_),
    .Q(execution_unit_0.register_file_0.r13_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09846_ (
    .CLK(dco_clk),
    .D(_01980_),
    .Q(execution_unit_0.register_file_0.r13_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09847_ (
    .CLK(dco_clk),
    .D(_01981_),
    .Q(execution_unit_0.register_file_0.r13_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09848_ (
    .CLK(dco_clk),
    .D(_01982_),
    .Q(execution_unit_0.register_file_0.r13_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09849_ (
    .CLK(dco_clk),
    .D(_01983_),
    .Q(execution_unit_0.register_file_0.r13_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09850_ (
    .CLK(dco_clk),
    .D(_01969_),
    .Q(execution_unit_0.register_file_0.r13_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09851_ (
    .CLK(dco_clk),
    .D(_01970_),
    .Q(execution_unit_0.register_file_0.r13_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09852_ (
    .CLK(dco_clk),
    .D(_01971_),
    .Q(execution_unit_0.register_file_0.r13_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09853_ (
    .CLK(dco_clk),
    .D(_01972_),
    .Q(execution_unit_0.register_file_0.r13_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09854_ (
    .CLK(dco_clk),
    .D(_01973_),
    .Q(execution_unit_0.register_file_0.r13_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09855_ (
    .CLK(dco_clk),
    .D(_01974_),
    .Q(execution_unit_0.register_file_0.r13_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09856_ (
    .CLK(dco_clk),
    .D(_01952_),
    .Q(execution_unit_0.register_file_0.r12_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09857_ (
    .CLK(dco_clk),
    .D(_01959_),
    .Q(execution_unit_0.register_file_0.r12_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09858_ (
    .CLK(dco_clk),
    .D(_01960_),
    .Q(execution_unit_0.register_file_0.r12_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09859_ (
    .CLK(dco_clk),
    .D(_01961_),
    .Q(execution_unit_0.register_file_0.r12_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09860_ (
    .CLK(dco_clk),
    .D(_01962_),
    .Q(execution_unit_0.register_file_0.r12_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09861_ (
    .CLK(dco_clk),
    .D(_01963_),
    .Q(execution_unit_0.register_file_0.r12_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09862_ (
    .CLK(dco_clk),
    .D(_01964_),
    .Q(execution_unit_0.register_file_0.r12_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09863_ (
    .CLK(dco_clk),
    .D(_01965_),
    .Q(execution_unit_0.register_file_0.r12_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09864_ (
    .CLK(dco_clk),
    .D(_01966_),
    .Q(execution_unit_0.register_file_0.r12_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09865_ (
    .CLK(dco_clk),
    .D(_01967_),
    .Q(execution_unit_0.register_file_0.r12_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09866_ (
    .CLK(dco_clk),
    .D(_01953_),
    .Q(execution_unit_0.register_file_0.r12_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09867_ (
    .CLK(dco_clk),
    .D(_01954_),
    .Q(execution_unit_0.register_file_0.r12_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09868_ (
    .CLK(dco_clk),
    .D(_01955_),
    .Q(execution_unit_0.register_file_0.r12_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09869_ (
    .CLK(dco_clk),
    .D(_01956_),
    .Q(execution_unit_0.register_file_0.r12_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09870_ (
    .CLK(dco_clk),
    .D(_01957_),
    .Q(execution_unit_0.register_file_0.r12_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09871_ (
    .CLK(dco_clk),
    .D(_01958_),
    .Q(execution_unit_0.register_file_0.r12_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09872_ (
    .CLK(dco_clk),
    .D(_01936_),
    .Q(execution_unit_0.register_file_0.r11_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09873_ (
    .CLK(dco_clk),
    .D(_01943_),
    .Q(execution_unit_0.register_file_0.r11_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09874_ (
    .CLK(dco_clk),
    .D(_01944_),
    .Q(execution_unit_0.register_file_0.r11_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09875_ (
    .CLK(dco_clk),
    .D(_01945_),
    .Q(execution_unit_0.register_file_0.r11_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09876_ (
    .CLK(dco_clk),
    .D(_01946_),
    .Q(execution_unit_0.register_file_0.r11_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09877_ (
    .CLK(dco_clk),
    .D(_01947_),
    .Q(execution_unit_0.register_file_0.r11_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09878_ (
    .CLK(dco_clk),
    .D(_01948_),
    .Q(execution_unit_0.register_file_0.r11_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09879_ (
    .CLK(dco_clk),
    .D(_01949_),
    .Q(execution_unit_0.register_file_0.r11_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09880_ (
    .CLK(dco_clk),
    .D(_01950_),
    .Q(execution_unit_0.register_file_0.r11_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09881_ (
    .CLK(dco_clk),
    .D(_01951_),
    .Q(execution_unit_0.register_file_0.r11_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09882_ (
    .CLK(dco_clk),
    .D(_01937_),
    .Q(execution_unit_0.register_file_0.r11_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09883_ (
    .CLK(dco_clk),
    .D(_01938_),
    .Q(execution_unit_0.register_file_0.r11_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09884_ (
    .CLK(dco_clk),
    .D(_01939_),
    .Q(execution_unit_0.register_file_0.r11_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09885_ (
    .CLK(dco_clk),
    .D(_01940_),
    .Q(execution_unit_0.register_file_0.r11_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09886_ (
    .CLK(dco_clk),
    .D(_01941_),
    .Q(execution_unit_0.register_file_0.r11_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09887_ (
    .CLK(dco_clk),
    .D(_01942_),
    .Q(execution_unit_0.register_file_0.r11_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09888_ (
    .CLK(dco_clk),
    .D(_01920_),
    .Q(execution_unit_0.register_file_0.r10_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09889_ (
    .CLK(dco_clk),
    .D(_01927_),
    .Q(execution_unit_0.register_file_0.r10_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09890_ (
    .CLK(dco_clk),
    .D(_01928_),
    .Q(execution_unit_0.register_file_0.r10_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09891_ (
    .CLK(dco_clk),
    .D(_01929_),
    .Q(execution_unit_0.register_file_0.r10_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09892_ (
    .CLK(dco_clk),
    .D(_01930_),
    .Q(execution_unit_0.register_file_0.r10_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09893_ (
    .CLK(dco_clk),
    .D(_01931_),
    .Q(execution_unit_0.register_file_0.r10_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09894_ (
    .CLK(dco_clk),
    .D(_01932_),
    .Q(execution_unit_0.register_file_0.r10_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09895_ (
    .CLK(dco_clk),
    .D(_01933_),
    .Q(execution_unit_0.register_file_0.r10_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09896_ (
    .CLK(dco_clk),
    .D(_01934_),
    .Q(execution_unit_0.register_file_0.r10_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09897_ (
    .CLK(dco_clk),
    .D(_01935_),
    .Q(execution_unit_0.register_file_0.r10_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09898_ (
    .CLK(dco_clk),
    .D(_01921_),
    .Q(execution_unit_0.register_file_0.r10_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09899_ (
    .CLK(dco_clk),
    .D(_01922_),
    .Q(execution_unit_0.register_file_0.r10_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09900_ (
    .CLK(dco_clk),
    .D(_01923_),
    .Q(execution_unit_0.register_file_0.r10_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09901_ (
    .CLK(dco_clk),
    .D(_01924_),
    .Q(execution_unit_0.register_file_0.r10_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09902_ (
    .CLK(dco_clk),
    .D(_01925_),
    .Q(execution_unit_0.register_file_0.r10_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09903_ (
    .CLK(dco_clk),
    .D(_01926_),
    .Q(execution_unit_0.register_file_0.r10_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09904_ (
    .CLK(dco_clk),
    .D(_02136_),
    .Q(execution_unit_0.register_file_0.r9_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09905_ (
    .CLK(dco_clk),
    .D(_02143_),
    .Q(execution_unit_0.register_file_0.r9_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09906_ (
    .CLK(dco_clk),
    .D(_02144_),
    .Q(execution_unit_0.register_file_0.r9_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09907_ (
    .CLK(dco_clk),
    .D(_02145_),
    .Q(execution_unit_0.register_file_0.r9_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09908_ (
    .CLK(dco_clk),
    .D(_02146_),
    .Q(execution_unit_0.register_file_0.r9_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09909_ (
    .CLK(dco_clk),
    .D(_02147_),
    .Q(execution_unit_0.register_file_0.r9_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09910_ (
    .CLK(dco_clk),
    .D(_02148_),
    .Q(execution_unit_0.register_file_0.r9_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09911_ (
    .CLK(dco_clk),
    .D(_02149_),
    .Q(execution_unit_0.register_file_0.r9_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09912_ (
    .CLK(dco_clk),
    .D(_02150_),
    .Q(execution_unit_0.register_file_0.r9_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09913_ (
    .CLK(dco_clk),
    .D(_02151_),
    .Q(execution_unit_0.register_file_0.r9_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09914_ (
    .CLK(dco_clk),
    .D(_02137_),
    .Q(execution_unit_0.register_file_0.r9_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09915_ (
    .CLK(dco_clk),
    .D(_02138_),
    .Q(execution_unit_0.register_file_0.r9_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09916_ (
    .CLK(dco_clk),
    .D(_02139_),
    .Q(execution_unit_0.register_file_0.r9_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09917_ (
    .CLK(dco_clk),
    .D(_02140_),
    .Q(execution_unit_0.register_file_0.r9_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09918_ (
    .CLK(dco_clk),
    .D(_02141_),
    .Q(execution_unit_0.register_file_0.r9_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09919_ (
    .CLK(dco_clk),
    .D(_02142_),
    .Q(execution_unit_0.register_file_0.r9_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09920_ (
    .CLK(dco_clk),
    .D(_02120_),
    .Q(execution_unit_0.register_file_0.r8_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09921_ (
    .CLK(dco_clk),
    .D(_02127_),
    .Q(execution_unit_0.register_file_0.r8_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09922_ (
    .CLK(dco_clk),
    .D(_02128_),
    .Q(execution_unit_0.register_file_0.r8_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09923_ (
    .CLK(dco_clk),
    .D(_02129_),
    .Q(execution_unit_0.register_file_0.r8_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09924_ (
    .CLK(dco_clk),
    .D(_02130_),
    .Q(execution_unit_0.register_file_0.r8_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09925_ (
    .CLK(dco_clk),
    .D(_02131_),
    .Q(execution_unit_0.register_file_0.r8_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09926_ (
    .CLK(dco_clk),
    .D(_02132_),
    .Q(execution_unit_0.register_file_0.r8_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09927_ (
    .CLK(dco_clk),
    .D(_02133_),
    .Q(execution_unit_0.register_file_0.r8_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09928_ (
    .CLK(dco_clk),
    .D(_02134_),
    .Q(execution_unit_0.register_file_0.r8_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09929_ (
    .CLK(dco_clk),
    .D(_02135_),
    .Q(execution_unit_0.register_file_0.r8_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09930_ (
    .CLK(dco_clk),
    .D(_02121_),
    .Q(execution_unit_0.register_file_0.r8_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09931_ (
    .CLK(dco_clk),
    .D(_02122_),
    .Q(execution_unit_0.register_file_0.r8_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09932_ (
    .CLK(dco_clk),
    .D(_02123_),
    .Q(execution_unit_0.register_file_0.r8_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09933_ (
    .CLK(dco_clk),
    .D(_02124_),
    .Q(execution_unit_0.register_file_0.r8_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09934_ (
    .CLK(dco_clk),
    .D(_02125_),
    .Q(execution_unit_0.register_file_0.r8_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09935_ (
    .CLK(dco_clk),
    .D(_02126_),
    .Q(execution_unit_0.register_file_0.r8_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09936_ (
    .CLK(dco_clk),
    .D(_02104_),
    .Q(execution_unit_0.register_file_0.r7_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09937_ (
    .CLK(dco_clk),
    .D(_02111_),
    .Q(execution_unit_0.register_file_0.r7_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09938_ (
    .CLK(dco_clk),
    .D(_02112_),
    .Q(execution_unit_0.register_file_0.r7_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09939_ (
    .CLK(dco_clk),
    .D(_02113_),
    .Q(execution_unit_0.register_file_0.r7_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09940_ (
    .CLK(dco_clk),
    .D(_02114_),
    .Q(execution_unit_0.register_file_0.r7_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09941_ (
    .CLK(dco_clk),
    .D(_02115_),
    .Q(execution_unit_0.register_file_0.r7_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09942_ (
    .CLK(dco_clk),
    .D(_02116_),
    .Q(execution_unit_0.register_file_0.r7_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09943_ (
    .CLK(dco_clk),
    .D(_02117_),
    .Q(execution_unit_0.register_file_0.r7_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09944_ (
    .CLK(dco_clk),
    .D(_02118_),
    .Q(execution_unit_0.register_file_0.r7_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09945_ (
    .CLK(dco_clk),
    .D(_02119_),
    .Q(execution_unit_0.register_file_0.r7_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09946_ (
    .CLK(dco_clk),
    .D(_02105_),
    .Q(execution_unit_0.register_file_0.r7_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09947_ (
    .CLK(dco_clk),
    .D(_02106_),
    .Q(execution_unit_0.register_file_0.r7_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09948_ (
    .CLK(dco_clk),
    .D(_02107_),
    .Q(execution_unit_0.register_file_0.r7_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09949_ (
    .CLK(dco_clk),
    .D(_02108_),
    .Q(execution_unit_0.register_file_0.r7_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09950_ (
    .CLK(dco_clk),
    .D(_02109_),
    .Q(execution_unit_0.register_file_0.r7_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09951_ (
    .CLK(dco_clk),
    .D(_02110_),
    .Q(execution_unit_0.register_file_0.r7_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09952_ (
    .CLK(dco_clk),
    .D(_02088_),
    .Q(execution_unit_0.register_file_0.r6_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09953_ (
    .CLK(dco_clk),
    .D(_02095_),
    .Q(execution_unit_0.register_file_0.r6_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09954_ (
    .CLK(dco_clk),
    .D(_02096_),
    .Q(execution_unit_0.register_file_0.r6_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09955_ (
    .CLK(dco_clk),
    .D(_02097_),
    .Q(execution_unit_0.register_file_0.r6_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09956_ (
    .CLK(dco_clk),
    .D(_02098_),
    .Q(execution_unit_0.register_file_0.r6_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09957_ (
    .CLK(dco_clk),
    .D(_02099_),
    .Q(execution_unit_0.register_file_0.r6_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09958_ (
    .CLK(dco_clk),
    .D(_02100_),
    .Q(execution_unit_0.register_file_0.r6_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09959_ (
    .CLK(dco_clk),
    .D(_02101_),
    .Q(execution_unit_0.register_file_0.r6_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09960_ (
    .CLK(dco_clk),
    .D(_02102_),
    .Q(execution_unit_0.register_file_0.r6_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09961_ (
    .CLK(dco_clk),
    .D(_02103_),
    .Q(execution_unit_0.register_file_0.r6_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09962_ (
    .CLK(dco_clk),
    .D(_02089_),
    .Q(execution_unit_0.register_file_0.r6_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09963_ (
    .CLK(dco_clk),
    .D(_02090_),
    .Q(execution_unit_0.register_file_0.r6_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09964_ (
    .CLK(dco_clk),
    .D(_02091_),
    .Q(execution_unit_0.register_file_0.r6_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09965_ (
    .CLK(dco_clk),
    .D(_02092_),
    .Q(execution_unit_0.register_file_0.r6_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09966_ (
    .CLK(dco_clk),
    .D(_02093_),
    .Q(execution_unit_0.register_file_0.r6_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09967_ (
    .CLK(dco_clk),
    .D(_02094_),
    .Q(execution_unit_0.register_file_0.r6_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09968_ (
    .CLK(dco_clk),
    .D(_02072_),
    .Q(execution_unit_0.register_file_0.r5_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09969_ (
    .CLK(dco_clk),
    .D(_02079_),
    .Q(execution_unit_0.register_file_0.r5_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09970_ (
    .CLK(dco_clk),
    .D(_02080_),
    .Q(execution_unit_0.register_file_0.r5_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09971_ (
    .CLK(dco_clk),
    .D(_02081_),
    .Q(execution_unit_0.register_file_0.r5_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09972_ (
    .CLK(dco_clk),
    .D(_02082_),
    .Q(execution_unit_0.register_file_0.r5_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09973_ (
    .CLK(dco_clk),
    .D(_02083_),
    .Q(execution_unit_0.register_file_0.r5_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09974_ (
    .CLK(dco_clk),
    .D(_02084_),
    .Q(execution_unit_0.register_file_0.r5_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09975_ (
    .CLK(dco_clk),
    .D(_02085_),
    .Q(execution_unit_0.register_file_0.r5_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09976_ (
    .CLK(dco_clk),
    .D(_02086_),
    .Q(execution_unit_0.register_file_0.r5_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09977_ (
    .CLK(dco_clk),
    .D(_02087_),
    .Q(execution_unit_0.register_file_0.r5_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09978_ (
    .CLK(dco_clk),
    .D(_02073_),
    .Q(execution_unit_0.register_file_0.r5_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09979_ (
    .CLK(dco_clk),
    .D(_02074_),
    .Q(execution_unit_0.register_file_0.r5_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09980_ (
    .CLK(dco_clk),
    .D(_02075_),
    .Q(execution_unit_0.register_file_0.r5_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09981_ (
    .CLK(dco_clk),
    .D(_02076_),
    .Q(execution_unit_0.register_file_0.r5_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09982_ (
    .CLK(dco_clk),
    .D(_02077_),
    .Q(execution_unit_0.register_file_0.r5_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09983_ (
    .CLK(dco_clk),
    .D(_02078_),
    .Q(execution_unit_0.register_file_0.r5_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09984_ (
    .CLK(dco_clk),
    .D(_02056_),
    .Q(execution_unit_0.register_file_0.r4_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09985_ (
    .CLK(dco_clk),
    .D(_02063_),
    .Q(execution_unit_0.register_file_0.r4_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09986_ (
    .CLK(dco_clk),
    .D(_02064_),
    .Q(execution_unit_0.register_file_0.r4_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09987_ (
    .CLK(dco_clk),
    .D(_02065_),
    .Q(execution_unit_0.register_file_0.r4_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09988_ (
    .CLK(dco_clk),
    .D(_02066_),
    .Q(execution_unit_0.register_file_0.r4_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09989_ (
    .CLK(dco_clk),
    .D(_02067_),
    .Q(execution_unit_0.register_file_0.r4_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09990_ (
    .CLK(dco_clk),
    .D(_02068_),
    .Q(execution_unit_0.register_file_0.r4_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09991_ (
    .CLK(dco_clk),
    .D(_02069_),
    .Q(execution_unit_0.register_file_0.r4_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09992_ (
    .CLK(dco_clk),
    .D(_02070_),
    .Q(execution_unit_0.register_file_0.r4_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09993_ (
    .CLK(dco_clk),
    .D(_02071_),
    .Q(execution_unit_0.register_file_0.r4_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09994_ (
    .CLK(dco_clk),
    .D(_02057_),
    .Q(execution_unit_0.register_file_0.r4_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09995_ (
    .CLK(dco_clk),
    .D(_02058_),
    .Q(execution_unit_0.register_file_0.r4_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09996_ (
    .CLK(dco_clk),
    .D(_02059_),
    .Q(execution_unit_0.register_file_0.r4_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09997_ (
    .CLK(dco_clk),
    .D(_02060_),
    .Q(execution_unit_0.register_file_0.r4_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09998_ (
    .CLK(dco_clk),
    .D(_02061_),
    .Q(execution_unit_0.register_file_0.r4_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _09999_ (
    .CLK(dco_clk),
    .D(_02062_),
    .Q(execution_unit_0.register_file_0.r4_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10000_ (
    .CLK(dco_clk),
    .D(_02040_),
    .Q(execution_unit_0.register_file_0.r3_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10001_ (
    .CLK(dco_clk),
    .D(_02047_),
    .Q(execution_unit_0.register_file_0.r3_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10002_ (
    .CLK(dco_clk),
    .D(_02048_),
    .Q(execution_unit_0.register_file_0.r3_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10003_ (
    .CLK(dco_clk),
    .D(_02049_),
    .Q(execution_unit_0.register_file_0.r3_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10004_ (
    .CLK(dco_clk),
    .D(_02050_),
    .Q(execution_unit_0.register_file_0.r3_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10005_ (
    .CLK(dco_clk),
    .D(_02051_),
    .Q(execution_unit_0.register_file_0.r3_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10006_ (
    .CLK(dco_clk),
    .D(_02052_),
    .Q(execution_unit_0.register_file_0.r3_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10007_ (
    .CLK(dco_clk),
    .D(_02053_),
    .Q(execution_unit_0.register_file_0.r3_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10008_ (
    .CLK(dco_clk),
    .D(_02054_),
    .Q(execution_unit_0.register_file_0.r3_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10009_ (
    .CLK(dco_clk),
    .D(_02055_),
    .Q(execution_unit_0.register_file_0.r3_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10010_ (
    .CLK(dco_clk),
    .D(_02041_),
    .Q(execution_unit_0.register_file_0.r3_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10011_ (
    .CLK(dco_clk),
    .D(_02042_),
    .Q(execution_unit_0.register_file_0.r3_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10012_ (
    .CLK(dco_clk),
    .D(_02043_),
    .Q(execution_unit_0.register_file_0.r3_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10013_ (
    .CLK(dco_clk),
    .D(_02044_),
    .Q(execution_unit_0.register_file_0.r3_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10014_ (
    .CLK(dco_clk),
    .D(_02045_),
    .Q(execution_unit_0.register_file_0.r3_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10015_ (
    .CLK(dco_clk),
    .D(_02046_),
    .Q(execution_unit_0.register_file_0.r3_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10016_ (
    .CLK(dco_clk),
    .D(_02032_),
    .Q(execution_unit_0.alu_0.status_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10017_ (
    .CLK(dco_clk),
    .D(_02033_),
    .Q(execution_unit_0.alu_0.status_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10018_ (
    .CLK(dco_clk),
    .D(_02034_),
    .Q(execution_unit_0.alu_0.status_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10019_ (
    .CLK(dco_clk),
    .D(_02035_),
    .Q(execution_unit_0.gie ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10020_ (
    .CLK(dco_clk),
    .D(_02036_),
    .Q(execution_unit_0.register_file_0.r2_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10021_ (
    .CLK(dco_clk),
    .D(_02037_),
    .Q(clock_module_0.oscoff ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10022_ (
    .CLK(dco_clk),
    .D(_02038_),
    .Q(clock_module_0.scg1 ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10023_ (
    .CLK(dco_clk),
    .D(_02039_),
    .Q(execution_unit_0.alu_0.status_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10024_ (
    .CLK(dco_clk),
    .D(_02016_),
    .Q(execution_unit_0.register_file_0.r1_0_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10025_ (
    .CLK(dco_clk),
    .D(_02023_),
    .Q(execution_unit_0.register_file_0.r1_1_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10026_ (
    .CLK(dco_clk),
    .D(_02024_),
    .Q(execution_unit_0.register_file_0.r1_2_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10027_ (
    .CLK(dco_clk),
    .D(_02025_),
    .Q(execution_unit_0.register_file_0.r1_3_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10028_ (
    .CLK(dco_clk),
    .D(_02026_),
    .Q(execution_unit_0.register_file_0.r1_4_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10029_ (
    .CLK(dco_clk),
    .D(_02027_),
    .Q(execution_unit_0.register_file_0.r1_5_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10030_ (
    .CLK(dco_clk),
    .D(_02028_),
    .Q(execution_unit_0.register_file_0.r1_6_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10031_ (
    .CLK(dco_clk),
    .D(_02029_),
    .Q(execution_unit_0.register_file_0.r1_7_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10032_ (
    .CLK(dco_clk),
    .D(_02030_),
    .Q(execution_unit_0.register_file_0.r1_8_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10033_ (
    .CLK(dco_clk),
    .D(_02031_),
    .Q(execution_unit_0.register_file_0.r1_9_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10034_ (
    .CLK(dco_clk),
    .D(_02017_),
    .Q(execution_unit_0.register_file_0.r1_10_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10035_ (
    .CLK(dco_clk),
    .D(_02018_),
    .Q(execution_unit_0.register_file_0.r1_11_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10036_ (
    .CLK(dco_clk),
    .D(_02019_),
    .Q(execution_unit_0.register_file_0.r1_12_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10037_ (
    .CLK(dco_clk),
    .D(_02020_),
    .Q(execution_unit_0.register_file_0.r1_13_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10038_ (
    .CLK(dco_clk),
    .D(_02021_),
    .Q(execution_unit_0.register_file_0.r1_14_ ),
    .R(_02152_),
    .S(1'h1)
  );
  DFFSR _10039_ (
    .CLK(dco_clk),
    .D(_02022_),
    .Q(execution_unit_0.register_file_0.r1_15_ ),
    .R(_02152_),
    .S(1'h1)
  );
  INVX1 _10040_ (
    .A(e_state_3_),
    .Y(_03624_)
  );
  INVX1 _10041_ (
    .A(e_state_2_),
    .Y(_03625_)
  );
  INVX1 _10042_ (
    .A(e_state_0_),
    .Y(_03626_)
  );
  INVX1 _10043_ (
    .A(execution_unit_0.gie ),
    .Y(_03627_)
  );
  INVX1 _10044_ (
    .A(irq_13_),
    .Y(_03628_)
  );
  INVX1 _10045_ (
    .A(irq_7_),
    .Y(_03629_)
  );
  INVX1 _10046_ (
    .A(irq_3_),
    .Y(_03630_)
  );
  INVX1 _10047_ (
    .A(irq_1_),
    .Y(_03631_)
  );
  INVX1 _10048_ (
    .A(cpu_halt_cmd),
    .Y(_03632_)
  );
  INVX1 _10049_ (
    .A(1'h0),
    .Y(_03633_)
  );
  INVX1 _10050_ (
    .A(frontend_0.i_state_4_ ),
    .Y(_03634_)
  );
  INVX1 _10051_ (
    .A(frontend_0.exec_dst_wr ),
    .Y(_03635_)
  );
  INVX1 _10052_ (
    .A(frontend_0.exec_jmp ),
    .Y(_03636_)
  );
  INVX1 _10053_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .Y(_03637_)
  );
  INVX1 _10054_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .Y(_03638_)
  );
  INVX1 _10055_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .Y(_03639_)
  );
  INVX1 _10056_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .Y(_03640_)
  );
  INVX1 _10057_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .Y(_03641_)
  );
  INVX1 _10058_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .Y(_03642_)
  );
  INVX1 _10059_ (
    .A(dbg_0.fe_mdb_in_0_ ),
    .Y(_03643_)
  );
  INVX1 _10060_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .Y(_03644_)
  );
  INVX1 _10061_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .Y(_03645_)
  );
  INVX1 _10062_ (
    .A(dbg_0.fe_mdb_in_3_ ),
    .Y(_03646_)
  );
  INVX1 _10063_ (
    .A(execution_unit_0.UNUSED_inst_ad_idx ),
    .Y(_03647_)
  );
  INVX1 _10064_ (
    .A(frontend_0.i_state_5_ ),
    .Y(_03648_)
  );
  INVX1 _10065_ (
    .A(frontend_0.i_state_2_ ),
    .Y(_03649_)
  );
  INVX1 _10066_ (
    .A(execution_unit_0.pc_sw_wr ),
    .Y(_03650_)
  );
  INVX1 _10067_ (
    .A(frontend_0.inst_sz_0_ ),
    .Y(_03651_)
  );
  INVX1 _10068_ (
    .A(frontend_0.i_state_1_ ),
    .Y(_03652_)
  );
  INVX1 _10069_ (
    .A(frontend_0.i_state_3_ ),
    .Y(_03653_)
  );
  INVX1 _10070_ (
    .A(frontend_0.i_state_0_ ),
    .Y(_03654_)
  );
  INVX1 _10071_ (
    .A(execution_unit_0.alu_0.alu_out_0_ ),
    .Y(_03655_)
  );
  INVX1 _10072_ (
    .A(dbg_0.UNUSED_pc_1_ ),
    .Y(_03656_)
  );
  INVX1 _10073_ (
    .A(frontend_0.irq_addr_1_ ),
    .Y(_03657_)
  );
  INVX1 _10074_ (
    .A(dbg_0.UNUSED_pc_2_ ),
    .Y(_03658_)
  );
  INVX1 _10075_ (
    .A(frontend_0.irq_addr_2_ ),
    .Y(_03659_)
  );
  INVX1 _10076_ (
    .A(dbg_0.UNUSED_pc_3_ ),
    .Y(_03660_)
  );
  INVX1 _10077_ (
    .A(frontend_0.irq_addr_3_ ),
    .Y(_03661_)
  );
  INVX1 _10078_ (
    .A(dbg_0.UNUSED_pc_4_ ),
    .Y(_03662_)
  );
  INVX1 _10079_ (
    .A(dbg_0.UNUSED_pc_5_ ),
    .Y(_03663_)
  );
  INVX1 _10080_ (
    .A(dbg_0.UNUSED_pc_6_ ),
    .Y(_03664_)
  );
  INVX1 _10081_ (
    .A(dbg_0.fe_mdb_in_6_ ),
    .Y(_03665_)
  );
  INVX1 _10082_ (
    .A(frontend_0.irq_addr_6_ ),
    .Y(_03666_)
  );
  INVX1 _10083_ (
    .A(dbg_0.UNUSED_pc_7_ ),
    .Y(_03667_)
  );
  INVX1 _10084_ (
    .A(dbg_0.UNUSED_pc_8_ ),
    .Y(_03668_)
  );
  INVX1 _10085_ (
    .A(dbg_0.UNUSED_pc_9_ ),
    .Y(_03669_)
  );
  INVX1 _10086_ (
    .A(dbg_0.UNUSED_pc_10_ ),
    .Y(_03670_)
  );
  INVX1 _10087_ (
    .A(dbg_0.UNUSED_pc_11_ ),
    .Y(_03671_)
  );
  INVX1 _10088_ (
    .A(dbg_0.UNUSED_pc_12_ ),
    .Y(_03672_)
  );
  INVX1 _10089_ (
    .A(dbg_0.fe_mdb_in_12_ ),
    .Y(_03673_)
  );
  INVX1 _10090_ (
    .A(dbg_0.UNUSED_pc_13_ ),
    .Y(_03674_)
  );
  INVX1 _10091_ (
    .A(dbg_0.UNUSED_pc_14_ ),
    .Y(_03675_)
  );
  INVX1 _10092_ (
    .A(dbg_0.UNUSED_pc_15_ ),
    .Y(_03676_)
  );
  INVX1 _10093_ (
    .A(frontend_0.inst_dest_bin_1_ ),
    .Y(_03677_)
  );
  INVX1 _10094_ (
    .A(frontend_0.inst_dest_bin_0_ ),
    .Y(_03678_)
  );
  INVX1 _10095_ (
    .A(frontend_0.inst_dest_bin_2_ ),
    .Y(_03679_)
  );
  INVX1 _10096_ (
    .A(frontend_0.inst_dest_bin_3_ ),
    .Y(_03680_)
  );
  INVX1 _10097_ (
    .A(execution_unit_0.inst_type_1_ ),
    .Y(_03681_)
  );
  INVX1 _10098_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .Y(_03682_)
  );
  INVX1 _10099_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .Y(_03683_)
  );
  INVX1 _10100_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .Y(_03684_)
  );
  INVX1 _10101_ (
    .A(dbg_0.dbg_mem_addr_2_ ),
    .Y(_03685_)
  );
  INVX1 _10102_ (
    .A(execution_unit_0.inst_type_0_ ),
    .Y(_03686_)
  );
  INVX1 _10103_ (
    .A(frontend_0.inst_src_bin_1_ ),
    .Y(_03687_)
  );
  INVX1 _10104_ (
    .A(frontend_0.inst_src_bin_3_ ),
    .Y(_03688_)
  );
  INVX1 _10105_ (
    .A(frontend_0.inst_src_bin_2_ ),
    .Y(_03689_)
  );
  INVX1 _10106_ (
    .A(execution_unit_0.inst_type_2_ ),
    .Y(_03690_)
  );
  INVX1 _10107_ (
    .A(execution_unit_0.alu_0.inst_alu_3_ ),
    .Y(_03691_)
  );
  INVX1 _10108_ (
    .A(execution_unit_0.alu_0.inst_alu_7_ ),
    .Y(_03692_)
  );
  INVX1 _10109_ (
    .A(execution_unit_0.alu_0.inst_alu_8_ ),
    .Y(_03693_)
  );
  INVX1 _10110_ (
    .A(frontend_0.inst_jmp_bin_0_ ),
    .Y(_03694_)
  );
  INVX1 _10111_ (
    .A(frontend_0.inst_jmp_bin_1_ ),
    .Y(_03695_)
  );
  INVX1 _10112_ (
    .A(execution_unit_0.inst_irq_rst ),
    .Y(_03696_)
  );
  INVX1 _10113_ (
    .A(_00162_),
    .Y(_03405_)
  );
  NOR2X1 _10114_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .Y(_03697_)
  );
  INVX1 _10115_ (
    .A(_03697_),
    .Y(_03698_)
  );
  NAND2X1 _10116_ (
    .A(e_state_3_),
    .B(e_state_2_),
    .Y(_03699_)
  );
  OAI21X1 _10117_ (
    .A(_03698_),
    .B(_03699_),
    .C(frontend_0.exec_jmp ),
    .Y(_03700_)
  );
  INVX1 _10118_ (
    .A(_03700_),
    .Y(_03701_)
  );
  NOR2X1 _10119_ (
    .A(_03624_),
    .B(e_state_2_),
    .Y(_03702_)
  );
  NAND2X1 _10120_ (
    .A(e_state_3_),
    .B(_03625_),
    .Y(_03703_)
  );
  NAND2X1 _10121_ (
    .A(_03626_),
    .B(e_state_1_),
    .Y(_03704_)
  );
  NOR2X1 _10122_ (
    .A(_03703_),
    .B(_03704_),
    .Y(_03705_)
  );
  OR2X1 _10123_ (
    .A(_03703_),
    .B(_03704_),
    .Y(_03706_)
  );
  OAI21X1 _10124_ (
    .A(_03703_),
    .B(_03704_),
    .C(frontend_0.exec_dst_wr ),
    .Y(_03707_)
  );
  AND2X1 _10125_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .Y(_03708_)
  );
  NAND2X1 _10126_ (
    .A(e_state_0_),
    .B(e_state_1_),
    .Y(_03709_)
  );
  NAND2X1 _10127_ (
    .A(_03624_),
    .B(e_state_2_),
    .Y(_03710_)
  );
  NOR2X1 _10128_ (
    .A(_03709_),
    .B(_03710_),
    .Y(_03711_)
  );
  NAND3X1 _10129_ (
    .A(_03624_),
    .B(e_state_2_),
    .C(_03708_),
    .Y(_03712_)
  );
  NAND3X1 _10130_ (
    .A(e_state_3_),
    .B(_03625_),
    .C(_03708_),
    .Y(_03713_)
  );
  MUX2X1 _10131_ (
    .A(_03712_),
    .B(_03713_),
    .S(frontend_0.exec_src_wr ),
    .Y(_03714_)
  );
  OAI21X1 _10132_ (
    .A(frontend_0.exec_dst_wr ),
    .B(_03714_),
    .C(_03707_),
    .Y(_03715_)
  );
  AOI21X1 _10133_ (
    .A(_03636_),
    .B(_03715_),
    .C(_03701_),
    .Y(exec_done)
  );
  NOR2X1 _10134_ (
    .A(frontend_0.i_state_4_ ),
    .B(exec_done),
    .Y(_03716_)
  );
  NOR2X1 _10135_ (
    .A(irq_12_),
    .B(irq_13_),
    .Y(_03717_)
  );
  NOR2X1 _10136_ (
    .A(irq_6_),
    .B(irq_7_),
    .Y(_03718_)
  );
  NOR2X1 _10137_ (
    .A(frontend_0.wdt_irq ),
    .B(irq_10_),
    .Y(_03719_)
  );
  NOR2X1 _10138_ (
    .A(irq_11_),
    .B(irq_9_),
    .Y(_03720_)
  );
  NAND2X1 _10139_ (
    .A(_03719_),
    .B(_03720_),
    .Y(_03721_)
  );
  NOR2X1 _10140_ (
    .A(irq_8_),
    .B(irq_2_),
    .Y(_03722_)
  );
  NAND3X1 _10141_ (
    .A(_03630_),
    .B(_03631_),
    .C(_03722_),
    .Y(_03723_)
  );
  NOR3X1 _10142_ (
    .A(irq_4_),
    .B(irq_5_),
    .C(irq_0_),
    .Y(_03724_)
  );
  NAND3X1 _10143_ (
    .A(_03717_),
    .B(_03718_),
    .C(_03724_),
    .Y(_03725_)
  );
  NOR3X1 _10144_ (
    .A(_03721_),
    .B(_03723_),
    .C(_03725_),
    .Y(_03726_)
  );
  OAI21X1 _10145_ (
    .A(_03627_),
    .B(_03726_),
    .C(_03633_),
    .Y(_03727_)
  );
  AND2X1 _10146_ (
    .A(cpu_en),
    .B(_03632_),
    .Y(_03728_)
  );
  NAND2X1 _10147_ (
    .A(cpu_en),
    .B(_03632_),
    .Y(_03729_)
  );
  NOR2X1 _10148_ (
    .A(cpu_halt_st),
    .B(_03729_),
    .Y(_03730_)
  );
  AND2X1 _10149_ (
    .A(_03727_),
    .B(_03730_),
    .Y(_03731_)
  );
  NAND2X1 _10150_ (
    .A(_03727_),
    .B(_03730_),
    .Y(_03732_)
  );
  NOR2X1 _10151_ (
    .A(_03716_),
    .B(_03732_),
    .Y(_03733_)
  );
  OAI21X1 _10152_ (
    .A(frontend_0.i_state_4_ ),
    .B(exec_done),
    .C(_03731_),
    .Y(_03734_)
  );
  NOR2X1 _10153_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(dbg_0.fe_mdb_in_14_ ),
    .Y(_03735_)
  );
  OAI21X1 _10154_ (
    .A(_03716_),
    .B(_03732_),
    .C(_03735_),
    .Y(_03736_)
  );
  NOR2X1 _10155_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_03736_),
    .Y(_03737_)
  );
  NAND3X1 _10156_ (
    .A(_03640_),
    .B(_03734_),
    .C(_03735_),
    .Y(_03738_)
  );
  NAND2X1 _10157_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(dbg_0.fe_mdb_in_7_ ),
    .Y(_03739_)
  );
  NOR2X1 _10158_ (
    .A(_03738_),
    .B(_03739_),
    .Y(_03740_)
  );
  OR2X1 _10159_ (
    .A(_03738_),
    .B(_03739_),
    .Y(_03741_)
  );
  AOI21X1 _10160_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03740_),
    .C(_03733_),
    .Y(_03742_)
  );
  NOR2X1 _10161_ (
    .A(cpu_halt_st),
    .B(_03742_),
    .Y(_03743_)
  );
  OR2X1 _10162_ (
    .A(cpu_halt_st),
    .B(_03742_),
    .Y(_03744_)
  );
  OR2X1 _10163_ (
    .A(_03640_),
    .B(_03736_),
    .Y(_03745_)
  );
  INVX1 _10164_ (
    .A(_03745_),
    .Y(_03746_)
  );
  AND2X1 _10165_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03745_),
    .Y(_03747_)
  );
  OAI21X1 _10166_ (
    .A(_03640_),
    .B(_03736_),
    .C(dbg_0.fe_mdb_in_5_ ),
    .Y(_03748_)
  );
  NAND2X1 _10167_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(_03747_),
    .Y(_03749_)
  );
  NOR2X1 _10168_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .B(dbg_0.fe_mdb_in_3_ ),
    .Y(_03750_)
  );
  NAND2X1 _10169_ (
    .A(_03645_),
    .B(_03646_),
    .Y(_03751_)
  );
  NOR2X1 _10170_ (
    .A(dbg_0.fe_mdb_in_10_ ),
    .B(dbg_0.fe_mdb_in_11_ ),
    .Y(_03752_)
  );
  INVX1 _10171_ (
    .A(_03752_),
    .Y(_03753_)
  );
  MUX2X1 _10172_ (
    .A(_03753_),
    .B(_03751_),
    .S(_03738_),
    .Y(_03754_)
  );
  MUX2X1 _10173_ (
    .A(_03752_),
    .B(_03750_),
    .S(_03738_),
    .Y(_03755_)
  );
  MUX2X1 _10174_ (
    .A(_03637_),
    .B(_03644_),
    .S(_03738_),
    .Y(_03756_)
  );
  MUX2X1 _10175_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(dbg_0.fe_mdb_in_1_ ),
    .S(_03738_),
    .Y(_03757_)
  );
  NOR2X1 _10176_ (
    .A(_03755_),
    .B(_03757_),
    .Y(_03758_)
  );
  NAND2X1 _10177_ (
    .A(_03754_),
    .B(_03756_),
    .Y(_03759_)
  );
  NOR2X1 _10178_ (
    .A(_03749_),
    .B(_03758_),
    .Y(_03760_)
  );
  NAND2X1 _10179_ (
    .A(_03642_),
    .B(_03747_),
    .Y(_03761_)
  );
  NAND2X1 _10180_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03639_),
    .Y(_03762_)
  );
  NOR2X1 _10181_ (
    .A(_03738_),
    .B(_03762_),
    .Y(_03763_)
  );
  INVX1 _10182_ (
    .A(_03763_),
    .Y(_03764_)
  );
  NAND2X1 _10183_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(_03763_),
    .Y(_03765_)
  );
  MUX2X1 _10184_ (
    .A(_03638_),
    .B(_03643_),
    .S(_03738_),
    .Y(_03766_)
  );
  MUX2X1 _10185_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(dbg_0.fe_mdb_in_0_ ),
    .S(_03738_),
    .Y(_03767_)
  );
  NAND3X1 _10186_ (
    .A(_03754_),
    .B(_03757_),
    .C(_03767_),
    .Y(_03768_)
  );
  NAND2X1 _10187_ (
    .A(_03760_),
    .B(_03768_),
    .Y(_03769_)
  );
  OR2X1 _10188_ (
    .A(_03749_),
    .B(_03768_),
    .Y(_03770_)
  );
  AOI22X1 _10189_ (
    .A(_03747_),
    .B(_03759_),
    .C(_03763_),
    .D(dbg_0.fe_mdb_in_8_ ),
    .Y(_03771_)
  );
  OAI21X1 _10190_ (
    .A(_03748_),
    .B(_03758_),
    .C(_03765_),
    .Y(_03772_)
  );
  NOR2X1 _10191_ (
    .A(_03733_),
    .B(_03735_),
    .Y(_03773_)
  );
  NAND2X1 _10192_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(_03773_),
    .Y(_03774_)
  );
  NOR2X1 _10193_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(_03738_),
    .Y(_03775_)
  );
  NAND2X1 _10194_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03775_),
    .Y(_03776_)
  );
  AOI21X1 _10195_ (
    .A(_03774_),
    .B(_03776_),
    .C(_03772_),
    .Y(_03777_)
  );
  OR2X1 _10196_ (
    .A(clock_module_0.UNUSED_cpuoff ),
    .B(_03729_),
    .Y(_03778_)
  );
  NOR2X1 _10197_ (
    .A(frontend_0.i_state_4_ ),
    .B(_03778_),
    .Y(_03779_)
  );
  OR2X1 _10198_ (
    .A(frontend_0.i_state_4_ ),
    .B(_03778_),
    .Y(_03780_)
  );
  NOR3X1 _10199_ (
    .A(_03755_),
    .B(_03757_),
    .C(_03767_),
    .Y(_03781_)
  );
  NAND3X1 _10200_ (
    .A(_03754_),
    .B(_03756_),
    .C(_03766_),
    .Y(_03782_)
  );
  OAI21X1 _10201_ (
    .A(_03640_),
    .B(_03736_),
    .C(dbg_0.fe_mdb_in_4_ ),
    .Y(_03783_)
  );
  NOR2X1 _10202_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03783_),
    .Y(_03784_)
  );
  OR2X1 _10203_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03783_),
    .Y(_03785_)
  );
  OAI21X1 _10204_ (
    .A(_03759_),
    .B(_03767_),
    .C(_03784_),
    .Y(_03786_)
  );
  AOI21X1 _10205_ (
    .A(_03782_),
    .B(_03784_),
    .C(_03780_),
    .Y(_03787_)
  );
  OAI21X1 _10206_ (
    .A(_03781_),
    .B(_03785_),
    .C(_03779_),
    .Y(_03788_)
  );
  OAI21X1 _10207_ (
    .A(_03777_),
    .B(_03788_),
    .C(_03744_),
    .Y(_03789_)
  );
  NOR2X1 _10208_ (
    .A(frontend_0.exec_jmp ),
    .B(_03713_),
    .Y(_03790_)
  );
  NOR2X1 _10209_ (
    .A(e_state_1_),
    .B(_03699_),
    .Y(_03791_)
  );
  NOR2X1 _10210_ (
    .A(_03711_),
    .B(_03791_),
    .Y(_03792_)
  );
  OAI21X1 _10211_ (
    .A(frontend_0.exec_jmp ),
    .B(_03706_),
    .C(_03792_),
    .Y(_03793_)
  );
  OAI21X1 _10212_ (
    .A(_03790_),
    .B(_03793_),
    .C(_03789_),
    .Y(_03794_)
  );
  OR2X1 _10213_ (
    .A(_03626_),
    .B(e_state_1_),
    .Y(_03795_)
  );
  NOR2X1 _10214_ (
    .A(_03703_),
    .B(_03795_),
    .Y(_03796_)
  );
  NOR2X1 _10215_ (
    .A(_03698_),
    .B(_03710_),
    .Y(_03797_)
  );
  NOR2X1 _10216_ (
    .A(_03796_),
    .B(_03797_),
    .Y(_03798_)
  );
  OAI21X1 _10217_ (
    .A(_03635_),
    .B(_03713_),
    .C(_03798_),
    .Y(_03799_)
  );
  NAND2X1 _10218_ (
    .A(_03624_),
    .B(_03625_),
    .Y(_03800_)
  );
  OR2X1 _10219_ (
    .A(e_state_0_),
    .B(_03800_),
    .Y(_03801_)
  );
  MUX2X1 _10220_ (
    .A(_03699_),
    .B(_03801_),
    .S(e_state_1_),
    .Y(_03802_)
  );
  NOR2X1 _10221_ (
    .A(_03799_),
    .B(_03802_),
    .Y(_03803_)
  );
  NOR2X1 _10222_ (
    .A(_03704_),
    .B(_03710_),
    .Y(_03804_)
  );
  NOR2X1 _10223_ (
    .A(execution_unit_0.UNUSED_inst_ad_symb ),
    .B(execution_unit_0.inst_ad_6_ ),
    .Y(_03805_)
  );
  NAND3X1 _10224_ (
    .A(_03647_),
    .B(_03804_),
    .C(_03805_),
    .Y(_03806_)
  );
  OR2X1 _10225_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .B(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .Y(_03807_)
  );
  OR2X1 _10226_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_03807_),
    .Y(_03808_)
  );
  NAND2X1 _10227_ (
    .A(frontend_0.exec_src_wr ),
    .B(_03790_),
    .Y(_03809_)
  );
  OAI21X1 _10228_ (
    .A(_03806_),
    .B(_03808_),
    .C(_03809_),
    .Y(_03810_)
  );
  NOR2X1 _10229_ (
    .A(execution_unit_0.inst_as_4_ ),
    .B(execution_unit_0.inst_as_1_ ),
    .Y(_03811_)
  );
  NOR2X1 _10230_ (
    .A(execution_unit_0.inst_as_6_ ),
    .B(execution_unit_0.inst_as_5_ ),
    .Y(_03812_)
  );
  NAND2X1 _10231_ (
    .A(_03811_),
    .B(_03812_),
    .Y(_03813_)
  );
  INVX1 _10232_ (
    .A(_03813_),
    .Y(_03814_)
  );
  NOR2X1 _10233_ (
    .A(_03648_),
    .B(_03814_),
    .Y(_03815_)
  );
  INVX1 _10234_ (
    .A(_03815_),
    .Y(_03816_)
  );
  OR2X1 _10235_ (
    .A(_03710_),
    .B(_03795_),
    .Y(_03817_)
  );
  INVX1 _10236_ (
    .A(_03817_),
    .Y(_03818_)
  );
  AOI21X1 _10237_ (
    .A(_03815_),
    .B(_03818_),
    .C(_03810_),
    .Y(_03819_)
  );
  NAND3X1 _10238_ (
    .A(_03794_),
    .B(_03803_),
    .C(_03819_),
    .Y(frontend_0.e_state_nxt_1_ )
  );
  OAI21X1 _10239_ (
    .A(frontend_0.i_state_4_ ),
    .B(frontend_0.i_state_2_ ),
    .C(_03733_),
    .Y(_03820_)
  );
  INVX1 _10240_ (
    .A(_03820_),
    .Y(_03402_)
  );
  NAND2X1 _10241_ (
    .A(e_state_0_),
    .B(_03791_),
    .Y(_03821_)
  );
  NOR2X1 _10242_ (
    .A(_03728_),
    .B(_03821_),
    .Y(_03822_)
  );
  OAI21X1 _10243_ (
    .A(exec_done),
    .B(_03822_),
    .C(_03778_),
    .Y(_03823_)
  );
  NAND3X1 _10244_ (
    .A(frontend_0.i_state_2_ ),
    .B(_03734_),
    .C(_03823_),
    .Y(_03824_)
  );
  AOI21X1 _10245_ (
    .A(_03648_),
    .B(_03824_),
    .C(_03650_),
    .Y(_03825_)
  );
  NAND3X1 _10246_ (
    .A(_03650_),
    .B(_03734_),
    .C(_03823_),
    .Y(_03826_)
  );
  INVX1 _10247_ (
    .A(_03826_),
    .Y(_03827_)
  );
  AOI21X1 _10248_ (
    .A(e_state_0_),
    .B(_03791_),
    .C(exec_done),
    .Y(_03828_)
  );
  NAND2X1 _10249_ (
    .A(frontend_0.i_state_2_ ),
    .B(_03828_),
    .Y(_03829_)
  );
  INVX1 _10250_ (
    .A(_03829_),
    .Y(_03830_)
  );
  NOR2X1 _10251_ (
    .A(_03634_),
    .B(_03778_),
    .Y(_03831_)
  );
  OR2X1 _10252_ (
    .A(_03651_),
    .B(frontend_0.inst_sz_1_ ),
    .Y(_03832_)
  );
  NOR2X1 _10253_ (
    .A(_03648_),
    .B(execution_unit_0.pc_sw_wr ),
    .Y(_03833_)
  );
  INVX1 _10254_ (
    .A(_03833_),
    .Y(_03834_)
  );
  NOR2X1 _10255_ (
    .A(frontend_0.i_state_1_ ),
    .B(frontend_0.i_state_3_ ),
    .Y(_03835_)
  );
  OAI21X1 _10256_ (
    .A(_03832_),
    .B(_03834_),
    .C(_03835_),
    .Y(_03836_)
  );
  AOI21X1 _10257_ (
    .A(_03732_),
    .B(_03831_),
    .C(_03836_),
    .Y(_03837_)
  );
  OAI21X1 _10258_ (
    .A(_03826_),
    .B(_03829_),
    .C(_03837_),
    .Y(_03838_)
  );
  NOR2X1 _10259_ (
    .A(_03825_),
    .B(_03838_),
    .Y(_03839_)
  );
  NOR2X1 _10260_ (
    .A(_03649_),
    .B(_03828_),
    .Y(dbg_0.decode_noirq )
  );
  NAND2X1 _10261_ (
    .A(_03827_),
    .B(dbg_0.decode_noirq ),
    .Y(_03840_)
  );
  NAND2X1 _10262_ (
    .A(_03839_),
    .B(_03840_),
    .Y(_03841_)
  );
  AND2X1 _10263_ (
    .A(_03770_),
    .B(_03786_),
    .Y(_03842_)
  );
  AND2X1 _10264_ (
    .A(_03774_),
    .B(_03842_),
    .Y(_03843_)
  );
  INVX1 _10265_ (
    .A(_03843_),
    .Y(_03844_)
  );
  OAI21X1 _10266_ (
    .A(_03840_),
    .B(_03844_),
    .C(_03839_),
    .Y(_03403_)
  );
  NAND2X1 _10267_ (
    .A(frontend_0.i_state_2_ ),
    .B(_03822_),
    .Y(_03845_)
  );
  OAI21X1 _10268_ (
    .A(frontend_0.i_state_4_ ),
    .B(frontend_0.i_state_2_ ),
    .C(_03778_),
    .Y(_03846_)
  );
  OR2X1 _10269_ (
    .A(_03731_),
    .B(_03846_),
    .Y(_03847_)
  );
  OAI21X1 _10270_ (
    .A(_03716_),
    .B(_03847_),
    .C(_03845_),
    .Y(_03404_)
  );
  NOR2X1 _10271_ (
    .A(_03840_),
    .B(_03843_),
    .Y(_03401_)
  );
  OAI21X1 _10272_ (
    .A(_03651_),
    .B(frontend_0.inst_sz_1_ ),
    .C(_03833_),
    .Y(_03848_)
  );
  INVX1 _10273_ (
    .A(_03848_),
    .Y(_03400_)
  );
  NAND2X1 _10274_ (
    .A(_03650_),
    .B(_03654_),
    .Y(_03849_)
  );
  AOI21X1 _10275_ (
    .A(_03643_),
    .B(frontend_0.i_state_3_ ),
    .C(_03849_),
    .Y(_03850_)
  );
  OAI21X1 _10276_ (
    .A(frontend_0.i_state_3_ ),
    .B(dbg_0.UNUSED_pc_0_ ),
    .C(_03850_),
    .Y(_03851_)
  );
  OAI21X1 _10277_ (
    .A(_03650_),
    .B(_03655_),
    .C(_03851_),
    .Y(UNUSED_fe_mab_0)
  );
  AOI21X1 _10278_ (
    .A(_03771_),
    .B(_03787_),
    .C(_03743_),
    .Y(_03852_)
  );
  OAI21X1 _10279_ (
    .A(_03772_),
    .B(_03788_),
    .C(_03744_),
    .Y(_03853_)
  );
  NOR3X1 _10280_ (
    .A(frontend_0.exec_src_wr ),
    .B(frontend_0.exec_jmp ),
    .C(_03852_),
    .Y(_03854_)
  );
  NOR2X1 _10281_ (
    .A(frontend_0.exec_dst_wr ),
    .B(_03713_),
    .Y(_03855_)
  );
  INVX1 _10282_ (
    .A(_03855_),
    .Y(_03856_)
  );
  NOR2X1 _10283_ (
    .A(_03854_),
    .B(_03856_),
    .Y(_03857_)
  );
  OR2X1 _10284_ (
    .A(_03854_),
    .B(_03856_),
    .Y(_03858_)
  );
  AOI21X1 _10285_ (
    .A(_03636_),
    .B(_03853_),
    .C(_03706_),
    .Y(_03859_)
  );
  NOR2X1 _10286_ (
    .A(_03709_),
    .B(_03800_),
    .Y(_03860_)
  );
  NOR2X1 _10287_ (
    .A(_03818_),
    .B(_03860_),
    .Y(_03861_)
  );
  OAI21X1 _10288_ (
    .A(_03792_),
    .B(_03853_),
    .C(_03861_),
    .Y(_03862_)
  );
  NOR2X1 _10289_ (
    .A(_03859_),
    .B(_03862_),
    .Y(_03863_)
  );
  OR2X1 _10290_ (
    .A(_03859_),
    .B(_03862_),
    .Y(_03864_)
  );
  OAI21X1 _10291_ (
    .A(_03854_),
    .B(_03856_),
    .C(_03863_),
    .Y(frontend_0.e_state_nxt_2_ )
  );
  NOR2X1 _10292_ (
    .A(_03650_),
    .B(execution_unit_0.alu_0.alu_out_1_ ),
    .Y(_03865_)
  );
  AOI21X1 _10293_ (
    .A(_03771_),
    .B(_03786_),
    .C(_03780_),
    .Y(_03866_)
  );
  OAI21X1 _10294_ (
    .A(frontend_0.exec_src_wr ),
    .B(_03713_),
    .C(_03792_),
    .Y(_03867_)
  );
  OAI21X1 _10295_ (
    .A(_03705_),
    .B(_03867_),
    .C(_03744_),
    .Y(_03868_)
  );
  NAND2X1 _10296_ (
    .A(e_state_1_),
    .B(frontend_0.exec_jmp ),
    .Y(_03869_)
  );
  NAND2X1 _10297_ (
    .A(_03697_),
    .B(_03702_),
    .Y(_03870_)
  );
  AOI21X1 _10298_ (
    .A(_03697_),
    .B(_03702_),
    .C(_03804_),
    .Y(_03871_)
  );
  OAI21X1 _10299_ (
    .A(_03703_),
    .B(_03869_),
    .C(_03871_),
    .Y(_03872_)
  );
  NOR2X1 _10300_ (
    .A(_03799_),
    .B(_03872_),
    .Y(_03873_)
  );
  OAI21X1 _10301_ (
    .A(_03866_),
    .B(_03868_),
    .C(_03873_),
    .Y(frontend_0.e_state_nxt_3_ )
  );
  AOI21X1 _10302_ (
    .A(_03771_),
    .B(_03774_),
    .C(_03788_),
    .Y(_03874_)
  );
  AND2X1 _10303_ (
    .A(_03635_),
    .B(_03790_),
    .Y(_03875_)
  );
  OAI21X1 _10304_ (
    .A(_03793_),
    .B(_03875_),
    .C(_03744_),
    .Y(_03876_)
  );
  AOI21X1 _10305_ (
    .A(frontend_0.i_state_5_ ),
    .B(_03814_),
    .C(frontend_0.i_state_1_ ),
    .Y(_03877_)
  );
  INVX1 _10306_ (
    .A(_03877_),
    .Y(_03878_)
  );
  NOR2X1 _10307_ (
    .A(frontend_0.exec_dext_rdy ),
    .B(_03878_),
    .Y(_03879_)
  );
  NOR2X1 _10308_ (
    .A(_03870_),
    .B(_03879_),
    .Y(_03880_)
  );
  NAND3X1 _10309_ (
    .A(_03798_),
    .B(_03801_),
    .C(_03806_),
    .Y(_03881_)
  );
  AOI21X1 _10310_ (
    .A(_03816_),
    .B(_03818_),
    .C(_03881_),
    .Y(_03882_)
  );
  OAI21X1 _10311_ (
    .A(frontend_0.exec_dst_wr ),
    .B(_03809_),
    .C(_03882_),
    .Y(_03883_)
  );
  NOR2X1 _10312_ (
    .A(_03880_),
    .B(_03883_),
    .Y(_03884_)
  );
  OAI21X1 _10313_ (
    .A(_03874_),
    .B(_03876_),
    .C(_03884_),
    .Y(frontend_0.e_state_nxt_0_ )
  );
  AND2X1 _10314_ (
    .A(frontend_0.e_state_nxt_3_ ),
    .B(frontend_0.e_state_nxt_0_ ),
    .Y(_03885_)
  );
  NAND2X1 _10315_ (
    .A(frontend_0.e_state_nxt_3_ ),
    .B(frontend_0.e_state_nxt_0_ ),
    .Y(_03886_)
  );
  AOI21X1 _10316_ (
    .A(_03858_),
    .B(_03863_),
    .C(_03886_),
    .Y(_03887_)
  );
  OAI21X1 _10317_ (
    .A(_03857_),
    .B(_03864_),
    .C(_03885_),
    .Y(_03888_)
  );
  OAI21X1 _10318_ (
    .A(_03830_),
    .B(_03887_),
    .C(_03656_),
    .Y(_03889_)
  );
  NOR3X1 _10319_ (
    .A(_03656_),
    .B(_03830_),
    .C(_03887_),
    .Y(_03890_)
  );
  NAND3X1 _10320_ (
    .A(dbg_0.UNUSED_pc_1_ ),
    .B(_03829_),
    .C(_03888_),
    .Y(_03891_)
  );
  AOI21X1 _10321_ (
    .A(_03889_),
    .B(_03891_),
    .C(frontend_0.i_state_3_ ),
    .Y(_03892_)
  );
  OAI21X1 _10322_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(_03653_),
    .C(_03654_),
    .Y(_03893_)
  );
  OR2X1 _10323_ (
    .A(_03892_),
    .B(_03893_),
    .Y(_03894_)
  );
  OAI21X1 _10324_ (
    .A(execution_unit_0.pc_sw_wr ),
    .B(frontend_0.irq_addr_1_ ),
    .C(_03849_),
    .Y(_03895_)
  );
  AOI21X1 _10325_ (
    .A(_03894_),
    .B(_03895_),
    .C(_03865_),
    .Y(execution_unit_0.pc_nxt_1_ )
  );
  NOR2X1 _10326_ (
    .A(_03650_),
    .B(execution_unit_0.alu_0.alu_out_2_ ),
    .Y(_03896_)
  );
  XNOR2X1 _10327_ (
    .A(_03658_),
    .B(_03890_),
    .Y(_03897_)
  );
  AOI21X1 _10328_ (
    .A(_03645_),
    .B(frontend_0.i_state_3_ ),
    .C(frontend_0.i_state_0_ ),
    .Y(_03898_)
  );
  OAI21X1 _10329_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03897_),
    .C(_03898_),
    .Y(_03899_)
  );
  AOI21X1 _10330_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_2_ ),
    .C(execution_unit_0.pc_sw_wr ),
    .Y(_03900_)
  );
  AOI21X1 _10331_ (
    .A(_03899_),
    .B(_03900_),
    .C(_03896_),
    .Y(execution_unit_0.pc_nxt_2_ )
  );
  OR2X1 _10332_ (
    .A(_03650_),
    .B(execution_unit_0.alu_0.alu_out_3_ ),
    .Y(_03901_)
  );
  OAI21X1 _10333_ (
    .A(_03658_),
    .B(_03891_),
    .C(_03660_),
    .Y(_03902_)
  );
  NOR3X1 _10334_ (
    .A(_03658_),
    .B(_03660_),
    .C(_03891_),
    .Y(_03903_)
  );
  NAND3X1 _10335_ (
    .A(dbg_0.UNUSED_pc_2_ ),
    .B(dbg_0.UNUSED_pc_3_ ),
    .C(_03890_),
    .Y(_03904_)
  );
  AOI21X1 _10336_ (
    .A(_03902_),
    .B(_03904_),
    .C(frontend_0.i_state_3_ ),
    .Y(_03905_)
  );
  OAI21X1 _10337_ (
    .A(dbg_0.fe_mdb_in_3_ ),
    .B(_03653_),
    .C(_03654_),
    .Y(_03906_)
  );
  OAI21X1 _10338_ (
    .A(execution_unit_0.pc_sw_wr ),
    .B(frontend_0.irq_addr_3_ ),
    .C(_03849_),
    .Y(_03907_)
  );
  OAI21X1 _10339_ (
    .A(_03905_),
    .B(_03906_),
    .C(_03907_),
    .Y(_03908_)
  );
  AND2X1 _10340_ (
    .A(_03901_),
    .B(_03908_),
    .Y(execution_unit_0.pc_nxt_3_ )
  );
  NOR2X1 _10341_ (
    .A(_03650_),
    .B(execution_unit_0.alu_0.alu_out_4_ ),
    .Y(_03909_)
  );
  XNOR2X1 _10342_ (
    .A(_03662_),
    .B(_03903_),
    .Y(_03910_)
  );
  AOI21X1 _10343_ (
    .A(_03642_),
    .B(frontend_0.i_state_3_ ),
    .C(frontend_0.i_state_0_ ),
    .Y(_03911_)
  );
  OAI21X1 _10344_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03910_),
    .C(_03911_),
    .Y(_03912_)
  );
  AOI21X1 _10345_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_4_ ),
    .C(execution_unit_0.pc_sw_wr ),
    .Y(_03913_)
  );
  AOI21X1 _10346_ (
    .A(_03912_),
    .B(_03913_),
    .C(_03909_),
    .Y(execution_unit_0.pc_nxt_4_ )
  );
  NOR2X1 _10347_ (
    .A(_03650_),
    .B(execution_unit_0.alu_0.alu_out_5_ ),
    .Y(_03914_)
  );
  NOR3X1 _10348_ (
    .A(_03662_),
    .B(_03663_),
    .C(_03904_),
    .Y(_03915_)
  );
  NAND3X1 _10349_ (
    .A(dbg_0.UNUSED_pc_4_ ),
    .B(dbg_0.UNUSED_pc_5_ ),
    .C(_03903_),
    .Y(_03916_)
  );
  OAI21X1 _10350_ (
    .A(_03662_),
    .B(_03904_),
    .C(_03663_),
    .Y(_03917_)
  );
  AOI21X1 _10351_ (
    .A(_03916_),
    .B(_03917_),
    .C(frontend_0.i_state_3_ ),
    .Y(_03918_)
  );
  OAI21X1 _10352_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03653_),
    .C(_03654_),
    .Y(_03919_)
  );
  OR2X1 _10353_ (
    .A(_03918_),
    .B(_03919_),
    .Y(_03920_)
  );
  NAND2X1 _10354_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_5_ ),
    .Y(_03921_)
  );
  AOI21X1 _10355_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_5_ ),
    .C(execution_unit_0.pc_sw_wr ),
    .Y(_03922_)
  );
  AOI21X1 _10356_ (
    .A(_03920_),
    .B(_03922_),
    .C(_03914_),
    .Y(execution_unit_0.pc_nxt_5_ )
  );
  NOR2X1 _10357_ (
    .A(_03650_),
    .B(execution_unit_0.alu_0.alu_out_6_ ),
    .Y(_03923_)
  );
  XNOR2X1 _10358_ (
    .A(_03664_),
    .B(_03915_),
    .Y(_03924_)
  );
  AOI21X1 _10359_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03665_),
    .C(frontend_0.i_state_0_ ),
    .Y(_03925_)
  );
  OAI21X1 _10360_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03924_),
    .C(_03925_),
    .Y(_03926_)
  );
  AOI21X1 _10361_ (
    .A(frontend_0.i_state_0_ ),
    .B(frontend_0.irq_addr_6_ ),
    .C(execution_unit_0.pc_sw_wr ),
    .Y(_03927_)
  );
  AOI21X1 _10362_ (
    .A(_03926_),
    .B(_03927_),
    .C(_03923_),
    .Y(execution_unit_0.pc_nxt_6_ )
  );
  NOR3X1 _10363_ (
    .A(_03664_),
    .B(_03667_),
    .C(_03916_),
    .Y(_03928_)
  );
  NAND3X1 _10364_ (
    .A(dbg_0.UNUSED_pc_6_ ),
    .B(dbg_0.UNUSED_pc_7_ ),
    .C(_03915_),
    .Y(_03929_)
  );
  OAI21X1 _10365_ (
    .A(_03664_),
    .B(_03916_),
    .C(_03667_),
    .Y(_03930_)
  );
  NAND2X1 _10366_ (
    .A(_03653_),
    .B(_03930_),
    .Y(_03931_)
  );
  AOI21X1 _10367_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03849_),
    .Y(_03932_)
  );
  OAI21X1 _10368_ (
    .A(_03928_),
    .B(_03931_),
    .C(_03932_),
    .Y(_03933_)
  );
  OAI21X1 _10369_ (
    .A(_03650_),
    .B(execution_unit_0.alu_0.alu_out_7_ ),
    .C(_03933_),
    .Y(_03934_)
  );
  INVX1 _10370_ (
    .A(_03934_),
    .Y(execution_unit_0.pc_nxt_7_ )
  );
  NOR2X1 _10371_ (
    .A(_03668_),
    .B(_03929_),
    .Y(_03935_)
  );
  OAI21X1 _10372_ (
    .A(dbg_0.UNUSED_pc_8_ ),
    .B(_03928_),
    .C(_03653_),
    .Y(_03936_)
  );
  AOI21X1 _10373_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03849_),
    .Y(_03937_)
  );
  OAI21X1 _10374_ (
    .A(_03935_),
    .B(_03936_),
    .C(_03937_),
    .Y(_03938_)
  );
  OAI21X1 _10375_ (
    .A(_03650_),
    .B(execution_unit_0.pc_sw_8_ ),
    .C(_03938_),
    .Y(_03939_)
  );
  INVX1 _10376_ (
    .A(_03939_),
    .Y(execution_unit_0.pc_nxt_8_ )
  );
  NOR3X1 _10377_ (
    .A(_03668_),
    .B(_03669_),
    .C(_03929_),
    .Y(_03940_)
  );
  NAND3X1 _10378_ (
    .A(dbg_0.UNUSED_pc_8_ ),
    .B(dbg_0.UNUSED_pc_9_ ),
    .C(_03928_),
    .Y(_03941_)
  );
  OAI21X1 _10379_ (
    .A(_03668_),
    .B(_03929_),
    .C(_03669_),
    .Y(_03942_)
  );
  NAND2X1 _10380_ (
    .A(_03653_),
    .B(_03942_),
    .Y(_03943_)
  );
  AOI21X1 _10381_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03849_),
    .Y(_03944_)
  );
  OAI21X1 _10382_ (
    .A(_03940_),
    .B(_03943_),
    .C(_03944_),
    .Y(_03945_)
  );
  OAI21X1 _10383_ (
    .A(_03650_),
    .B(execution_unit_0.pc_sw_9_ ),
    .C(_03945_),
    .Y(_03946_)
  );
  INVX1 _10384_ (
    .A(_03946_),
    .Y(execution_unit_0.pc_nxt_9_ )
  );
  XNOR2X1 _10385_ (
    .A(dbg_0.UNUSED_pc_10_ ),
    .B(_03940_),
    .Y(_03947_)
  );
  AOI21X1 _10386_ (
    .A(dbg_0.fe_mdb_in_10_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03849_),
    .Y(_03948_)
  );
  OAI21X1 _10387_ (
    .A(frontend_0.i_state_3_ ),
    .B(_03947_),
    .C(_03948_),
    .Y(_03949_)
  );
  OAI21X1 _10388_ (
    .A(_03650_),
    .B(execution_unit_0.pc_sw_10_ ),
    .C(_03949_),
    .Y(_03950_)
  );
  INVX1 _10389_ (
    .A(_03950_),
    .Y(execution_unit_0.pc_nxt_10_ )
  );
  NOR3X1 _10390_ (
    .A(_03670_),
    .B(_03671_),
    .C(_03941_),
    .Y(_03951_)
  );
  NAND3X1 _10391_ (
    .A(dbg_0.UNUSED_pc_10_ ),
    .B(dbg_0.UNUSED_pc_11_ ),
    .C(_03940_),
    .Y(_03952_)
  );
  OAI21X1 _10392_ (
    .A(_03670_),
    .B(_03941_),
    .C(_03671_),
    .Y(_03953_)
  );
  NAND2X1 _10393_ (
    .A(_03653_),
    .B(_03953_),
    .Y(_03954_)
  );
  AOI21X1 _10394_ (
    .A(dbg_0.fe_mdb_in_11_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03849_),
    .Y(_03955_)
  );
  OAI21X1 _10395_ (
    .A(_03951_),
    .B(_03954_),
    .C(_03955_),
    .Y(_03956_)
  );
  OAI21X1 _10396_ (
    .A(_03650_),
    .B(execution_unit_0.pc_sw_11_ ),
    .C(_03956_),
    .Y(_03957_)
  );
  INVX1 _10397_ (
    .A(_03957_),
    .Y(execution_unit_0.pc_nxt_11_ )
  );
  NOR2X1 _10398_ (
    .A(_03650_),
    .B(execution_unit_0.pc_sw_12_ ),
    .Y(_03958_)
  );
  AOI21X1 _10399_ (
    .A(_03672_),
    .B(_03952_),
    .C(frontend_0.i_state_3_ ),
    .Y(_03959_)
  );
  OAI21X1 _10400_ (
    .A(_03672_),
    .B(_03952_),
    .C(_03959_),
    .Y(_03960_)
  );
  AOI21X1 _10401_ (
    .A(frontend_0.i_state_3_ ),
    .B(dbg_0.fe_mdb_in_12_ ),
    .C(_03849_),
    .Y(_03961_)
  );
  AOI21X1 _10402_ (
    .A(_03960_),
    .B(_03961_),
    .C(_03958_),
    .Y(execution_unit_0.pc_nxt_12_ )
  );
  NOR2X1 _10403_ (
    .A(_03650_),
    .B(execution_unit_0.pc_sw_13_ ),
    .Y(_03962_)
  );
  NOR3X1 _10404_ (
    .A(_03672_),
    .B(_03674_),
    .C(_03952_),
    .Y(_03963_)
  );
  NAND3X1 _10405_ (
    .A(dbg_0.UNUSED_pc_12_ ),
    .B(dbg_0.UNUSED_pc_13_ ),
    .C(_03951_),
    .Y(_03964_)
  );
  OAI21X1 _10406_ (
    .A(_03672_),
    .B(_03952_),
    .C(_03674_),
    .Y(_03965_)
  );
  NAND3X1 _10407_ (
    .A(_03653_),
    .B(_03964_),
    .C(_03965_),
    .Y(_03966_)
  );
  AOI21X1 _10408_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03849_),
    .Y(_03967_)
  );
  AOI21X1 _10409_ (
    .A(_03966_),
    .B(_03967_),
    .C(_03962_),
    .Y(execution_unit_0.pc_nxt_13_ )
  );
  NOR2X1 _10410_ (
    .A(_03650_),
    .B(execution_unit_0.pc_sw_14_ ),
    .Y(_03968_)
  );
  AOI21X1 _10411_ (
    .A(_03675_),
    .B(_03964_),
    .C(frontend_0.i_state_3_ ),
    .Y(_03969_)
  );
  OAI21X1 _10412_ (
    .A(_03675_),
    .B(_03964_),
    .C(_03969_),
    .Y(_03970_)
  );
  AOI21X1 _10413_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03849_),
    .Y(_03971_)
  );
  AOI21X1 _10414_ (
    .A(_03970_),
    .B(_03971_),
    .C(_03968_),
    .Y(execution_unit_0.pc_nxt_14_ )
  );
  NOR2X1 _10415_ (
    .A(_03650_),
    .B(execution_unit_0.pc_sw_15_ ),
    .Y(_03972_)
  );
  OAI21X1 _10416_ (
    .A(_03675_),
    .B(_03964_),
    .C(_03676_),
    .Y(_03973_)
  );
  NAND3X1 _10417_ (
    .A(dbg_0.UNUSED_pc_14_ ),
    .B(dbg_0.UNUSED_pc_15_ ),
    .C(_03963_),
    .Y(_03974_)
  );
  NAND3X1 _10418_ (
    .A(_03653_),
    .B(_03973_),
    .C(_03974_),
    .Y(_03975_)
  );
  AOI21X1 _10419_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(frontend_0.i_state_3_ ),
    .C(_03849_),
    .Y(_03976_)
  );
  AOI21X1 _10420_ (
    .A(_03975_),
    .B(_03976_),
    .C(_03972_),
    .Y(execution_unit_0.pc_nxt_15_ )
  );
  NOR2X1 _10421_ (
    .A(frontend_0.inst_dest_bin_2_ ),
    .B(frontend_0.inst_dest_bin_3_ ),
    .Y(_03977_)
  );
  NOR2X1 _10422_ (
    .A(frontend_0.inst_dest_bin_1_ ),
    .B(frontend_0.inst_dest_bin_0_ ),
    .Y(_03978_)
  );
  AND2X1 _10423_ (
    .A(_03977_),
    .B(_03978_),
    .Y(_03979_)
  );
  NOR2X1 _10424_ (
    .A(execution_unit_0.alu_0.inst_so_7_ ),
    .B(_03807_),
    .Y(_03980_)
  );
  INVX1 _10425_ (
    .A(_03980_),
    .Y(_03981_)
  );
  AOI21X1 _10426_ (
    .A(_03979_),
    .B(_03980_),
    .C(execution_unit_0.inst_type_1_ ),
    .Y(_03982_)
  );
  NAND2X1 _10427_ (
    .A(_03682_),
    .B(_03683_),
    .Y(_03983_)
  );
  NAND3X1 _10428_ (
    .A(cpu_halt_st),
    .B(_03684_),
    .C(_03685_),
    .Y(_03984_)
  );
  OAI22X1 _10429_ (
    .A(cpu_halt_st),
    .B(_03982_),
    .C(_03983_),
    .D(_03984_),
    .Y(execution_unit_0.inst_dest_0_ )
  );
  NOR2X1 _10430_ (
    .A(frontend_0.inst_dest_bin_1_ ),
    .B(_03678_),
    .Y(_03985_)
  );
  AND2X1 _10431_ (
    .A(_03977_),
    .B(_03985_),
    .Y(_03986_)
  );
  NOR2X1 _10432_ (
    .A(cpu_halt_st),
    .B(execution_unit_0.inst_type_1_ ),
    .Y(_03987_)
  );
  OAI21X1 _10433_ (
    .A(_03981_),
    .B(_03986_),
    .C(_03987_),
    .Y(_03988_)
  );
  NAND2X1 _10434_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .B(_03683_),
    .Y(_03989_)
  );
  OAI21X1 _10435_ (
    .A(_03984_),
    .B(_03989_),
    .C(_03988_),
    .Y(execution_unit_0.inst_dest_1_ )
  );
  NOR2X1 _10436_ (
    .A(_03677_),
    .B(frontend_0.inst_dest_bin_0_ ),
    .Y(_03990_)
  );
  NAND2X1 _10437_ (
    .A(_03977_),
    .B(_03990_),
    .Y(_03991_)
  );
  NAND2X1 _10438_ (
    .A(_03980_),
    .B(_03987_),
    .Y(_03992_)
  );
  NAND2X1 _10439_ (
    .A(_03682_),
    .B(dbg_0.dbg_mem_addr_1_ ),
    .Y(_03993_)
  );
  OAI22X1 _10440_ (
    .A(_03991_),
    .B(_03992_),
    .C(_03993_),
    .D(_03984_),
    .Y(execution_unit_0.inst_dest_2_ )
  );
  NOR2X1 _10441_ (
    .A(_03677_),
    .B(_03678_),
    .Y(_03994_)
  );
  NAND2X1 _10442_ (
    .A(_03977_),
    .B(_03994_),
    .Y(_03995_)
  );
  NAND2X1 _10443_ (
    .A(dbg_0.dbg_mem_addr_0_ ),
    .B(dbg_0.dbg_mem_addr_1_ ),
    .Y(_03996_)
  );
  OAI22X1 _10444_ (
    .A(_03992_),
    .B(_03995_),
    .C(_03996_),
    .D(_03984_),
    .Y(execution_unit_0.inst_dest_3_ )
  );
  NOR2X1 _10445_ (
    .A(_03679_),
    .B(frontend_0.inst_dest_bin_3_ ),
    .Y(_03997_)
  );
  NAND2X1 _10446_ (
    .A(_03978_),
    .B(_03997_),
    .Y(_03998_)
  );
  NAND2X1 _10447_ (
    .A(_03684_),
    .B(dbg_0.dbg_mem_addr_2_ ),
    .Y(_03999_)
  );
  NAND3X1 _10448_ (
    .A(cpu_halt_st),
    .B(_03682_),
    .C(_03683_),
    .Y(_04000_)
  );
  OAI22X1 _10449_ (
    .A(_03992_),
    .B(_03998_),
    .C(_03999_),
    .D(_04000_),
    .Y(execution_unit_0.inst_dest_4_ )
  );
  NAND2X1 _10450_ (
    .A(_03985_),
    .B(_03997_),
    .Y(_04001_)
  );
  NAND3X1 _10451_ (
    .A(cpu_halt_st),
    .B(dbg_0.dbg_mem_addr_0_ ),
    .C(_03683_),
    .Y(_04002_)
  );
  OAI22X1 _10452_ (
    .A(_03992_),
    .B(_04001_),
    .C(_04002_),
    .D(_03999_),
    .Y(execution_unit_0.inst_dest_5_ )
  );
  NAND2X1 _10453_ (
    .A(_03990_),
    .B(_03997_),
    .Y(_04003_)
  );
  NAND3X1 _10454_ (
    .A(cpu_halt_st),
    .B(_03682_),
    .C(dbg_0.dbg_mem_addr_1_ ),
    .Y(_04004_)
  );
  OAI22X1 _10455_ (
    .A(_03992_),
    .B(_04003_),
    .C(_04004_),
    .D(_03999_),
    .Y(execution_unit_0.inst_dest_6_ )
  );
  NAND2X1 _10456_ (
    .A(_03994_),
    .B(_03997_),
    .Y(_04005_)
  );
  NAND3X1 _10457_ (
    .A(cpu_halt_st),
    .B(dbg_0.dbg_mem_addr_0_ ),
    .C(dbg_0.dbg_mem_addr_1_ ),
    .Y(_04006_)
  );
  OAI22X1 _10458_ (
    .A(_03992_),
    .B(_04005_),
    .C(_04006_),
    .D(_03999_),
    .Y(execution_unit_0.inst_dest_7_ )
  );
  NOR2X1 _10459_ (
    .A(frontend_0.inst_dest_bin_2_ ),
    .B(_03680_),
    .Y(_04007_)
  );
  NAND2X1 _10460_ (
    .A(_03978_),
    .B(_04007_),
    .Y(_04008_)
  );
  NAND2X1 _10461_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .B(_03685_),
    .Y(_04009_)
  );
  OAI22X1 _10462_ (
    .A(_03992_),
    .B(_04008_),
    .C(_04009_),
    .D(_04000_),
    .Y(execution_unit_0.inst_dest_8_ )
  );
  NAND2X1 _10463_ (
    .A(_03985_),
    .B(_04007_),
    .Y(_04010_)
  );
  OAI22X1 _10464_ (
    .A(_04002_),
    .B(_04009_),
    .C(_04010_),
    .D(_03992_),
    .Y(execution_unit_0.inst_dest_9_ )
  );
  NAND2X1 _10465_ (
    .A(_03990_),
    .B(_04007_),
    .Y(_04011_)
  );
  OAI22X1 _10466_ (
    .A(_04004_),
    .B(_04009_),
    .C(_04011_),
    .D(_03992_),
    .Y(execution_unit_0.inst_dest_10_ )
  );
  NAND2X1 _10467_ (
    .A(_03994_),
    .B(_04007_),
    .Y(_04012_)
  );
  OAI22X1 _10468_ (
    .A(_04006_),
    .B(_04009_),
    .C(_04012_),
    .D(_03992_),
    .Y(execution_unit_0.inst_dest_11_ )
  );
  NOR2X1 _10469_ (
    .A(_03679_),
    .B(_03680_),
    .Y(_04013_)
  );
  NAND2X1 _10470_ (
    .A(_03978_),
    .B(_04013_),
    .Y(_04014_)
  );
  NAND2X1 _10471_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .B(dbg_0.dbg_mem_addr_2_ ),
    .Y(_04015_)
  );
  OAI22X1 _10472_ (
    .A(_03992_),
    .B(_04014_),
    .C(_04015_),
    .D(_04000_),
    .Y(execution_unit_0.inst_dest_12_ )
  );
  NAND2X1 _10473_ (
    .A(_03985_),
    .B(_04013_),
    .Y(_04016_)
  );
  OAI22X1 _10474_ (
    .A(_04002_),
    .B(_04015_),
    .C(_04016_),
    .D(_03992_),
    .Y(execution_unit_0.inst_dest_13_ )
  );
  NAND2X1 _10475_ (
    .A(_03990_),
    .B(_04013_),
    .Y(_04017_)
  );
  OAI22X1 _10476_ (
    .A(_04004_),
    .B(_04015_),
    .C(_04017_),
    .D(_03992_),
    .Y(execution_unit_0.inst_dest_14_ )
  );
  NAND2X1 _10477_ (
    .A(_03994_),
    .B(_04013_),
    .Y(_04018_)
  );
  OAI22X1 _10478_ (
    .A(_04006_),
    .B(_04015_),
    .C(_04018_),
    .D(_03992_),
    .Y(execution_unit_0.inst_dest_15_ )
  );
  AND2X1 _10479_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(_03979_),
    .Y(_04019_)
  );
  NOR2X1 _10480_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(execution_unit_0.inst_type_2_ ),
    .Y(_04020_)
  );
  OAI21X1 _10481_ (
    .A(execution_unit_0.alu_0.inst_so_7_ ),
    .B(_04019_),
    .C(_04020_),
    .Y(_04021_)
  );
  OR2X1 _10482_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(frontend_0.inst_src_bin_1_ ),
    .Y(_04022_)
  );
  NAND3X1 _10483_ (
    .A(_03688_),
    .B(_03689_),
    .C(execution_unit_0.inst_type_2_ ),
    .Y(_04023_)
  );
  OAI21X1 _10484_ (
    .A(_04022_),
    .B(_04023_),
    .C(_04021_),
    .Y(execution_unit_0.inst_src_0_ )
  );
  NOR2X1 _10485_ (
    .A(execution_unit_0.alu_0.inst_so_7_ ),
    .B(_03686_),
    .Y(_04024_)
  );
  AOI21X1 _10486_ (
    .A(_03986_),
    .B(_04024_),
    .C(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .Y(_04025_)
  );
  NAND2X1 _10487_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(_03687_),
    .Y(_04026_)
  );
  OAI22X1 _10488_ (
    .A(execution_unit_0.inst_type_2_ ),
    .B(_04025_),
    .C(_04026_),
    .D(_04023_),
    .Y(execution_unit_0.inst_src_1_ )
  );
  NAND2X1 _10489_ (
    .A(_04020_),
    .B(_04024_),
    .Y(_04027_)
  );
  OR2X1 _10490_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(_03687_),
    .Y(_04028_)
  );
  OAI22X1 _10491_ (
    .A(_03991_),
    .B(_04027_),
    .C(_04028_),
    .D(_04023_),
    .Y(execution_unit_0.inst_src_2_ )
  );
  NAND2X1 _10492_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(frontend_0.inst_src_bin_1_ ),
    .Y(_04029_)
  );
  OAI22X1 _10493_ (
    .A(_03995_),
    .B(_04027_),
    .C(_04029_),
    .D(_04023_),
    .Y(execution_unit_0.inst_src_3_ )
  );
  NAND2X1 _10494_ (
    .A(_03688_),
    .B(frontend_0.inst_src_bin_2_ ),
    .Y(_04030_)
  );
  OR2X1 _10495_ (
    .A(_03690_),
    .B(_04022_),
    .Y(_04031_)
  );
  OAI22X1 _10496_ (
    .A(_03998_),
    .B(_04027_),
    .C(_04030_),
    .D(_04031_),
    .Y(execution_unit_0.inst_src_4_ )
  );
  OR2X1 _10497_ (
    .A(_03690_),
    .B(_04026_),
    .Y(_04032_)
  );
  OAI22X1 _10498_ (
    .A(_04001_),
    .B(_04027_),
    .C(_04030_),
    .D(_04032_),
    .Y(execution_unit_0.inst_src_5_ )
  );
  OR2X1 _10499_ (
    .A(_03690_),
    .B(_04028_),
    .Y(_04033_)
  );
  OAI22X1 _10500_ (
    .A(_04003_),
    .B(_04027_),
    .C(_04030_),
    .D(_04033_),
    .Y(execution_unit_0.inst_src_6_ )
  );
  OR2X1 _10501_ (
    .A(_03690_),
    .B(_04029_),
    .Y(_04034_)
  );
  OAI22X1 _10502_ (
    .A(_04005_),
    .B(_04027_),
    .C(_04030_),
    .D(_04034_),
    .Y(execution_unit_0.inst_src_7_ )
  );
  NAND2X1 _10503_ (
    .A(frontend_0.inst_src_bin_3_ ),
    .B(_03689_),
    .Y(_04035_)
  );
  OAI22X1 _10504_ (
    .A(_04008_),
    .B(_04027_),
    .C(_04031_),
    .D(_04035_),
    .Y(execution_unit_0.inst_src_8_ )
  );
  OAI22X1 _10505_ (
    .A(_04010_),
    .B(_04027_),
    .C(_04032_),
    .D(_04035_),
    .Y(execution_unit_0.inst_src_9_ )
  );
  OAI22X1 _10506_ (
    .A(_04011_),
    .B(_04027_),
    .C(_04033_),
    .D(_04035_),
    .Y(execution_unit_0.inst_src_10_ )
  );
  OAI22X1 _10507_ (
    .A(_04012_),
    .B(_04027_),
    .C(_04034_),
    .D(_04035_),
    .Y(execution_unit_0.inst_src_11_ )
  );
  NAND2X1 _10508_ (
    .A(frontend_0.inst_src_bin_3_ ),
    .B(frontend_0.inst_src_bin_2_ ),
    .Y(_04036_)
  );
  OAI22X1 _10509_ (
    .A(_04014_),
    .B(_04027_),
    .C(_04031_),
    .D(_04036_),
    .Y(execution_unit_0.inst_src_12_ )
  );
  OAI22X1 _10510_ (
    .A(_04016_),
    .B(_04027_),
    .C(_04032_),
    .D(_04036_),
    .Y(execution_unit_0.inst_src_13_ )
  );
  OAI22X1 _10511_ (
    .A(_04017_),
    .B(_04027_),
    .C(_04033_),
    .D(_04036_),
    .Y(execution_unit_0.inst_src_14_ )
  );
  OAI22X1 _10512_ (
    .A(_04018_),
    .B(_04027_),
    .C(_04034_),
    .D(_04036_),
    .Y(execution_unit_0.inst_src_15_ )
  );
  NOR2X1 _10513_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .Y(_04037_)
  );
  OAI21X1 _10514_ (
    .A(_03649_),
    .B(_03828_),
    .C(_03734_),
    .Y(_04038_)
  );
  AND2X1 _10515_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03734_),
    .Y(_04039_)
  );
  OAI21X1 _10516_ (
    .A(_03716_),
    .B(_03732_),
    .C(dbg_0.fe_mdb_in_15_ ),
    .Y(_04040_)
  );
  NAND2X1 _10517_ (
    .A(_03641_),
    .B(_04039_),
    .Y(_04041_)
  );
  NOR2X1 _10518_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(dbg_0.fe_mdb_in_12_ ),
    .Y(_04042_)
  );
  OAI21X1 _10519_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_04041_),
    .C(_04038_),
    .Y(_04043_)
  );
  NAND2X1 _10520_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(dbg_0.fe_mdb_in_12_ ),
    .Y(_04044_)
  );
  NOR2X1 _10521_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03641_),
    .Y(_04045_)
  );
  AND2X1 _10522_ (
    .A(_03734_),
    .B(_04045_),
    .Y(_04046_)
  );
  INVX1 _10523_ (
    .A(_04046_),
    .Y(_04047_)
  );
  NAND2X1 _10524_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .B(_04039_),
    .Y(_04048_)
  );
  NAND3X1 _10525_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .B(_04039_),
    .C(_04042_),
    .Y(_04049_)
  );
  OAI21X1 _10526_ (
    .A(_04044_),
    .B(_04047_),
    .C(_04049_),
    .Y(_04050_)
  );
  OAI22X1 _10527_ (
    .A(execution_unit_0.alu_0.inst_alu_0_ ),
    .B(_04038_),
    .C(_04043_),
    .D(_04050_),
    .Y(_04051_)
  );
  INVX1 _10528_ (
    .A(_04051_),
    .Y(_03316_)
  );
  OAI21X1 _10529_ (
    .A(execution_unit_0.alu_0.inst_alu_1_ ),
    .B(_04038_),
    .C(_04043_),
    .Y(_04052_)
  );
  INVX1 _10530_ (
    .A(_04052_),
    .Y(_03319_)
  );
  NAND2X1 _10531_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(dbg_0.decode_noirq ),
    .Y(_04053_)
  );
  OR2X1 _10532_ (
    .A(dbg_0.fe_mdb_in_12_ ),
    .B(_04053_),
    .Y(_04054_)
  );
  OR2X1 _10533_ (
    .A(_04041_),
    .B(_04054_),
    .Y(_04055_)
  );
  OAI21X1 _10534_ (
    .A(_04047_),
    .B(_04053_),
    .C(_04055_),
    .Y(_04056_)
  );
  AOI21X1 _10535_ (
    .A(execution_unit_0.alu_0.inst_alu_2_ ),
    .B(_04037_),
    .C(_04056_),
    .Y(_04057_)
  );
  INVX1 _10536_ (
    .A(_04057_),
    .Y(_03320_)
  );
  OAI21X1 _10537_ (
    .A(_03640_),
    .B(_03736_),
    .C(_03765_),
    .Y(_04058_)
  );
  OAI22X1 _10538_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_04041_),
    .C(_04042_),
    .D(_04047_),
    .Y(_04059_)
  );
  OAI21X1 _10539_ (
    .A(_04058_),
    .B(_04059_),
    .C(_04038_),
    .Y(_04060_)
  );
  OAI21X1 _10540_ (
    .A(_03691_),
    .B(_04038_),
    .C(_04060_),
    .Y(_03321_)
  );
  NOR2X1 _10541_ (
    .A(execution_unit_0.alu_0.inst_alu_4_ ),
    .B(_04038_),
    .Y(_04061_)
  );
  NOR2X1 _10542_ (
    .A(_04040_),
    .B(_04044_),
    .Y(_04062_)
  );
  NOR2X1 _10543_ (
    .A(_04037_),
    .B(_04062_),
    .Y(_04063_)
  );
  AOI21X1 _10544_ (
    .A(_04049_),
    .B(_04063_),
    .C(_04061_),
    .Y(_03322_)
  );
  NAND2X1 _10545_ (
    .A(execution_unit_0.alu_0.inst_alu_5_ ),
    .B(_04037_),
    .Y(_04064_)
  );
  NAND2X1 _10546_ (
    .A(_03773_),
    .B(dbg_0.decode_noirq ),
    .Y(_04065_)
  );
  NOR2X1 _10547_ (
    .A(_03641_),
    .B(_03673_),
    .Y(_04066_)
  );
  NAND3X1 _10548_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03640_),
    .C(_04066_),
    .Y(_04067_)
  );
  OAI21X1 _10549_ (
    .A(_04065_),
    .B(_04067_),
    .C(_04064_),
    .Y(_03323_)
  );
  NAND2X1 _10550_ (
    .A(execution_unit_0.alu_0.inst_alu_6_ ),
    .B(_04037_),
    .Y(_04068_)
  );
  OAI21X1 _10551_ (
    .A(_04048_),
    .B(_04054_),
    .C(_04068_),
    .Y(_03324_)
  );
  OAI21X1 _10552_ (
    .A(_03692_),
    .B(_04038_),
    .C(_04055_),
    .Y(_03325_)
  );
  NOR2X1 _10553_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03741_),
    .Y(_04069_)
  );
  OAI21X1 _10554_ (
    .A(_04062_),
    .B(_04069_),
    .C(_04038_),
    .Y(_04070_)
  );
  OAI21X1 _10555_ (
    .A(_03693_),
    .B(_04038_),
    .C(_04070_),
    .Y(_03326_)
  );
  NOR2X1 _10556_ (
    .A(execution_unit_0.alu_0.inst_alu_9_ ),
    .B(_04038_),
    .Y(_04071_)
  );
  AOI21X1 _10557_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_04039_),
    .C(_04059_),
    .Y(_04072_)
  );
  NOR2X1 _10558_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(dbg_0.fe_mdb_in_7_ ),
    .Y(_04073_)
  );
  INVX1 _10559_ (
    .A(_04073_),
    .Y(_04074_)
  );
  AOI21X1 _10560_ (
    .A(_03737_),
    .B(_04073_),
    .C(_04037_),
    .Y(_04075_)
  );
  OAI21X1 _10561_ (
    .A(_03738_),
    .B(_04074_),
    .C(_04038_),
    .Y(_04076_)
  );
  NOR2X1 _10562_ (
    .A(_04069_),
    .B(_04076_),
    .Y(_04077_)
  );
  AOI21X1 _10563_ (
    .A(_04072_),
    .B(_04077_),
    .C(_04071_),
    .Y(_03327_)
  );
  OAI21X1 _10564_ (
    .A(execution_unit_0.alu_0.inst_alu_10_ ),
    .B(_04038_),
    .C(_04076_),
    .Y(_04078_)
  );
  INVX1 _10565_ (
    .A(_04078_),
    .Y(_03317_)
  );
  NAND2X1 _10566_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_alu ),
    .B(_04037_),
    .Y(_04079_)
  );
  NAND3X1 _10567_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03641_),
    .C(dbg_0.fe_mdb_in_12_ ),
    .Y(_04080_)
  );
  OAI21X1 _10568_ (
    .A(_04065_),
    .B(_04080_),
    .C(_04079_),
    .Y(_03318_)
  );
  NOR2X1 _10569_ (
    .A(_03796_),
    .B(_03879_),
    .Y(_03308_)
  );
  NAND2X1 _10570_ (
    .A(execution_unit_0.inst_ad_0_ ),
    .B(_04037_),
    .Y(_04081_)
  );
  OAI21X1 _10571_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(_04065_),
    .C(_04081_),
    .Y(_03312_)
  );
  OR2X1 _10572_ (
    .A(_03639_),
    .B(_04065_),
    .Y(_04082_)
  );
  NOR2X1 _10573_ (
    .A(dbg_0.fe_mdb_in_0_ ),
    .B(_03751_),
    .Y(_04083_)
  );
  OAI22X1 _10574_ (
    .A(_03647_),
    .B(_04038_),
    .C(_04082_),
    .D(_04083_),
    .Y(_03313_)
  );
  NAND2X1 _10575_ (
    .A(execution_unit_0.UNUSED_inst_ad_symb ),
    .B(_04037_),
    .Y(_04084_)
  );
  NAND2X1 _10576_ (
    .A(_03644_),
    .B(_04083_),
    .Y(_04085_)
  );
  OAI21X1 _10577_ (
    .A(_04082_),
    .B(_04085_),
    .C(_04084_),
    .Y(_03314_)
  );
  NAND2X1 _10578_ (
    .A(execution_unit_0.inst_ad_6_ ),
    .B(_04037_),
    .Y(_04086_)
  );
  NAND2X1 _10579_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(_04083_),
    .Y(_04087_)
  );
  OAI21X1 _10580_ (
    .A(_04082_),
    .B(_04087_),
    .C(_04086_),
    .Y(_03315_)
  );
  OAI21X1 _10581_ (
    .A(_03774_),
    .B(_03842_),
    .C(_04038_),
    .Y(_04088_)
  );
  OAI22X1 _10582_ (
    .A(_03651_),
    .B(_04038_),
    .C(_04088_),
    .D(_03843_),
    .Y(_03389_)
  );
  OAI21X1 _10583_ (
    .A(frontend_0.inst_sz_1_ ),
    .B(_04038_),
    .C(_04088_),
    .Y(_04089_)
  );
  INVX1 _10584_ (
    .A(_04089_),
    .Y(_03390_)
  );
  NAND2X1 _10585_ (
    .A(execution_unit_0.alu_0.inst_bw ),
    .B(_04037_),
    .Y(_04090_)
  );
  NOR2X1 _10586_ (
    .A(_03665_),
    .B(_03733_),
    .Y(_04091_)
  );
  NAND3X1 _10587_ (
    .A(_03745_),
    .B(dbg_0.decode_noirq ),
    .C(_04091_),
    .Y(_04092_)
  );
  OAI21X1 _10588_ (
    .A(_03729_),
    .B(_04092_),
    .C(_04090_),
    .Y(_03336_)
  );
  NOR2X1 _10589_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(dbg_0.fe_mdb_in_5_ ),
    .Y(_04093_)
  );
  NOR2X1 _10590_ (
    .A(execution_unit_0.inst_as_0_ ),
    .B(_04038_),
    .Y(_04094_)
  );
  AOI21X1 _10591_ (
    .A(_03782_),
    .B(_04093_),
    .C(_04037_),
    .Y(_04095_)
  );
  AOI21X1 _10592_ (
    .A(_03745_),
    .B(_04095_),
    .C(_04094_),
    .Y(_03328_)
  );
  OAI21X1 _10593_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .C(_03784_),
    .Y(_04096_)
  );
  NOR2X1 _10594_ (
    .A(_03758_),
    .B(_04096_),
    .Y(_04097_)
  );
  AOI22X1 _10595_ (
    .A(execution_unit_0.inst_as_1_ ),
    .B(_04037_),
    .C(_04097_),
    .D(_03768_),
    .Y(_04098_)
  );
  INVX1 _10596_ (
    .A(_04098_),
    .Y(_03329_)
  );
  OAI21X1 _10597_ (
    .A(_03758_),
    .B(_03761_),
    .C(_04038_),
    .Y(_04099_)
  );
  OAI21X1 _10598_ (
    .A(execution_unit_0.inst_as_2_ ),
    .B(_04038_),
    .C(_04099_),
    .Y(_04100_)
  );
  INVX1 _10599_ (
    .A(_04100_),
    .Y(_03330_)
  );
  NAND2X1 _10600_ (
    .A(execution_unit_0.inst_as_3_ ),
    .B(_04037_),
    .Y(_04101_)
  );
  OAI21X1 _10601_ (
    .A(_03769_),
    .B(_04037_),
    .C(_04101_),
    .Y(_03331_)
  );
  NAND2X1 _10602_ (
    .A(execution_unit_0.inst_as_4_ ),
    .B(_04037_),
    .Y(_04102_)
  );
  OAI21X1 _10603_ (
    .A(_03768_),
    .B(_04096_),
    .C(_04102_),
    .Y(_03332_)
  );
  NAND2X1 _10604_ (
    .A(execution_unit_0.inst_as_5_ ),
    .B(_04037_),
    .Y(_04103_)
  );
  OAI21X1 _10605_ (
    .A(_03770_),
    .B(_04037_),
    .C(_04103_),
    .Y(_03333_)
  );
  NAND2X1 _10606_ (
    .A(_03758_),
    .B(_03767_),
    .Y(_04104_)
  );
  NAND2X1 _10607_ (
    .A(execution_unit_0.inst_as_6_ ),
    .B(_04037_),
    .Y(_04105_)
  );
  OAI21X1 _10608_ (
    .A(_04096_),
    .B(_04104_),
    .C(_04105_),
    .Y(_03334_)
  );
  OAI21X1 _10609_ (
    .A(_03640_),
    .B(_03736_),
    .C(_03781_),
    .Y(_04106_)
  );
  OAI21X1 _10610_ (
    .A(_03748_),
    .B(_04104_),
    .C(_04106_),
    .Y(_04107_)
  );
  AND2X1 _10611_ (
    .A(_04038_),
    .B(_04107_),
    .Y(_04108_)
  );
  AOI21X1 _10612_ (
    .A(execution_unit_0.inst_as_7_ ),
    .B(_04037_),
    .C(_04108_),
    .Y(_04109_)
  );
  INVX1 _10613_ (
    .A(_04109_),
    .Y(_03335_)
  );
  NAND2X1 _10614_ (
    .A(execution_unit_0.inst_mov ),
    .B(_04037_),
    .Y(_04110_)
  );
  NAND2X1 _10615_ (
    .A(_04042_),
    .B(_04045_),
    .Y(_04111_)
  );
  OAI21X1 _10616_ (
    .A(_04065_),
    .B(_04111_),
    .C(_04110_),
    .Y(_03361_)
  );
  OAI21X1 _10617_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .C(_03638_),
    .Y(_04112_)
  );
  OAI21X1 _10618_ (
    .A(frontend_0.inst_src_bin_0_ ),
    .B(_04038_),
    .C(_04112_),
    .Y(_04113_)
  );
  INVX1 _10619_ (
    .A(_04113_),
    .Y(_03385_)
  );
  OAI21X1 _10620_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .C(_03637_),
    .Y(_04114_)
  );
  OAI21X1 _10621_ (
    .A(frontend_0.inst_src_bin_1_ ),
    .B(_04038_),
    .C(_04114_),
    .Y(_04115_)
  );
  INVX1 _10622_ (
    .A(_04115_),
    .Y(_03386_)
  );
  OAI21X1 _10623_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_10_ ),
    .Y(_04116_)
  );
  OAI21X1 _10624_ (
    .A(_03689_),
    .B(_04038_),
    .C(_04116_),
    .Y(_03387_)
  );
  OAI21X1 _10625_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_11_ ),
    .Y(_04117_)
  );
  OAI21X1 _10626_ (
    .A(_03688_),
    .B(_04038_),
    .C(_04117_),
    .Y(_03388_)
  );
  OAI21X1 _10627_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_0_ ),
    .Y(_04118_)
  );
  OAI21X1 _10628_ (
    .A(_03678_),
    .B(_04038_),
    .C(_04118_),
    .Y(_03337_)
  );
  OAI21X1 _10629_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_1_ ),
    .Y(_04119_)
  );
  OAI21X1 _10630_ (
    .A(_03677_),
    .B(_04038_),
    .C(_04119_),
    .Y(_03338_)
  );
  OAI21X1 _10631_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_2_ ),
    .Y(_04120_)
  );
  OAI21X1 _10632_ (
    .A(_03679_),
    .B(_04038_),
    .C(_04120_),
    .Y(_03339_)
  );
  OAI21X1 _10633_ (
    .A(_03733_),
    .B(dbg_0.decode_noirq ),
    .C(dbg_0.fe_mdb_in_3_ ),
    .Y(_04121_)
  );
  OAI21X1 _10634_ (
    .A(_03680_),
    .B(_04038_),
    .C(_04121_),
    .Y(_03340_)
  );
  NAND2X1 _10635_ (
    .A(_03737_),
    .B(dbg_0.decode_noirq ),
    .Y(_04122_)
  );
  OAI21X1 _10636_ (
    .A(_03686_),
    .B(_04038_),
    .C(_04122_),
    .Y(_03391_)
  );
  AND2X1 _10637_ (
    .A(_03746_),
    .B(dbg_0.decode_noirq ),
    .Y(_04123_)
  );
  NAND2X1 _10638_ (
    .A(_03746_),
    .B(dbg_0.decode_noirq ),
    .Y(_04124_)
  );
  OAI21X1 _10639_ (
    .A(_03681_),
    .B(_04038_),
    .C(_04124_),
    .Y(_03392_)
  );
  OAI21X1 _10640_ (
    .A(_03690_),
    .B(_04038_),
    .C(_04065_),
    .Y(_03393_)
  );
  OAI21X1 _10641_ (
    .A(_03694_),
    .B(_04038_),
    .C(_04116_),
    .Y(_03358_)
  );
  OAI21X1 _10642_ (
    .A(_03695_),
    .B(_04038_),
    .C(_04117_),
    .Y(_03359_)
  );
  NAND2X1 _10643_ (
    .A(frontend_0.inst_jmp_bin_2_ ),
    .B(_04037_),
    .Y(_04125_)
  );
  OAI21X1 _10644_ (
    .A(_03673_),
    .B(_04037_),
    .C(_04125_),
    .Y(_03360_)
  );
  NAND2X1 _10645_ (
    .A(execution_unit_0.alu_0.inst_so_0_ ),
    .B(_04037_),
    .Y(_04126_)
  );
  AOI21X1 _10646_ (
    .A(_04112_),
    .B(_04126_),
    .C(_04075_),
    .Y(_03378_)
  );
  NAND2X1 _10647_ (
    .A(execution_unit_0.alu_0.inst_so_1_ ),
    .B(_04037_),
    .Y(_04127_)
  );
  NAND3X1 _10648_ (
    .A(_03637_),
    .B(_03775_),
    .C(_04038_),
    .Y(_04128_)
  );
  OAI21X1 _10649_ (
    .A(_03639_),
    .B(_04128_),
    .C(_04127_),
    .Y(_03379_)
  );
  NAND2X1 _10650_ (
    .A(execution_unit_0.alu_0.inst_so_3_ ),
    .B(_04037_),
    .Y(_04129_)
  );
  OAI21X1 _10651_ (
    .A(_03741_),
    .B(_04114_),
    .C(_04129_),
    .Y(_03380_)
  );
  NAND2X1 _10652_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .B(_04037_),
    .Y(_04130_)
  );
  OAI21X1 _10653_ (
    .A(_03764_),
    .B(_04112_),
    .C(_04130_),
    .Y(_03381_)
  );
  NAND3X1 _10654_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03638_),
    .C(dbg_0.fe_mdb_in_7_ ),
    .Y(_04131_)
  );
  NAND2X1 _10655_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .B(_04037_),
    .Y(_04132_)
  );
  OAI21X1 _10656_ (
    .A(_04122_),
    .B(_04131_),
    .C(_04132_),
    .Y(_03382_)
  );
  NAND2X1 _10657_ (
    .A(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .B(_04037_),
    .Y(_04133_)
  );
  OAI21X1 _10658_ (
    .A(_03765_),
    .B(_04037_),
    .C(_04133_),
    .Y(_03383_)
  );
  NOR2X1 _10659_ (
    .A(execution_unit_0.alu_0.inst_so_7_ ),
    .B(_04038_),
    .Y(_04134_)
  );
  AOI21X1 _10660_ (
    .A(_03742_),
    .B(_04038_),
    .C(_04134_),
    .Y(_03384_)
  );
  MUX2X1 _10661_ (
    .A(execution_unit_0.inst_dext_0_ ),
    .B(dbg_0.fe_mdb_in_0_ ),
    .S(_03877_),
    .Y(_04135_)
  );
  INVX1 _10662_ (
    .A(_04135_),
    .Y(_03341_)
  );
  NAND2X1 _10663_ (
    .A(execution_unit_0.inst_dext_1_ ),
    .B(_03877_),
    .Y(_04136_)
  );
  NOR2X1 _10664_ (
    .A(frontend_0.i_state_0_ ),
    .B(_03404_),
    .Y(_04137_)
  );
  OAI21X1 _10665_ (
    .A(_03840_),
    .B(_03843_),
    .C(_04137_),
    .Y(_04138_)
  );
  NAND3X1 _10666_ (
    .A(_03839_),
    .B(_03840_),
    .C(_04137_),
    .Y(_04139_)
  );
  OAI21X1 _10667_ (
    .A(_03848_),
    .B(_04139_),
    .C(frontend_0.i_state_5_ ),
    .Y(_04140_)
  );
  OAI21X1 _10668_ (
    .A(execution_unit_0.inst_as_4_ ),
    .B(_04140_),
    .C(_03652_),
    .Y(_03406_)
  );
  AOI22X1 _10669_ (
    .A(frontend_0.i_state_5_ ),
    .B(execution_unit_0.inst_as_4_ ),
    .C(_03406_),
    .D(execution_unit_0.UNUSED_inst_ad_symb ),
    .Y(_03407_)
  );
  OR2X1 _10670_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(_03407_),
    .Y(_03408_)
  );
  XNOR2X1 _10671_ (
    .A(_03644_),
    .B(_03407_),
    .Y(_03409_)
  );
  OAI21X1 _10672_ (
    .A(_03877_),
    .B(_03409_),
    .C(_04136_),
    .Y(_03348_)
  );
  NAND2X1 _10673_ (
    .A(execution_unit_0.inst_dext_2_ ),
    .B(_03877_),
    .Y(_03410_)
  );
  NOR2X1 _10674_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .B(_03408_),
    .Y(_03411_)
  );
  XNOR2X1 _10675_ (
    .A(_03645_),
    .B(_03408_),
    .Y(_03412_)
  );
  OAI21X1 _10676_ (
    .A(_03877_),
    .B(_03412_),
    .C(_03410_),
    .Y(_03349_)
  );
  OAI21X1 _10677_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .B(_03408_),
    .C(dbg_0.fe_mdb_in_3_ ),
    .Y(_03413_)
  );
  NAND2X1 _10678_ (
    .A(_03646_),
    .B(_03411_),
    .Y(_03414_)
  );
  AND2X1 _10679_ (
    .A(_03413_),
    .B(_03414_),
    .Y(_03415_)
  );
  NAND2X1 _10680_ (
    .A(execution_unit_0.inst_dext_3_ ),
    .B(_03877_),
    .Y(_03416_)
  );
  OAI21X1 _10681_ (
    .A(_03877_),
    .B(_03415_),
    .C(_03416_),
    .Y(_03350_)
  );
  NAND2X1 _10682_ (
    .A(execution_unit_0.inst_dext_4_ ),
    .B(_03877_),
    .Y(_03417_)
  );
  XNOR2X1 _10683_ (
    .A(_03642_),
    .B(_03414_),
    .Y(_03418_)
  );
  OAI21X1 _10684_ (
    .A(_03877_),
    .B(_03418_),
    .C(_03417_),
    .Y(_03351_)
  );
  OAI21X1 _10685_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(_03414_),
    .C(dbg_0.fe_mdb_in_5_ ),
    .Y(_03419_)
  );
  NAND3X1 _10686_ (
    .A(_03646_),
    .B(_04093_),
    .C(_03411_),
    .Y(_03420_)
  );
  AND2X1 _10687_ (
    .A(_03419_),
    .B(_03420_),
    .Y(_03421_)
  );
  NAND2X1 _10688_ (
    .A(execution_unit_0.inst_dext_5_ ),
    .B(_03877_),
    .Y(_03422_)
  );
  OAI21X1 _10689_ (
    .A(_03877_),
    .B(_03421_),
    .C(_03422_),
    .Y(_03352_)
  );
  NAND2X1 _10690_ (
    .A(execution_unit_0.inst_dext_6_ ),
    .B(_03877_),
    .Y(_03423_)
  );
  NOR2X1 _10691_ (
    .A(dbg_0.fe_mdb_in_6_ ),
    .B(_03420_),
    .Y(_03424_)
  );
  XNOR2X1 _10692_ (
    .A(_03665_),
    .B(_03420_),
    .Y(_03425_)
  );
  OAI21X1 _10693_ (
    .A(_03877_),
    .B(_03425_),
    .C(_03423_),
    .Y(_03353_)
  );
  OAI21X1 _10694_ (
    .A(dbg_0.fe_mdb_in_6_ ),
    .B(_03420_),
    .C(dbg_0.fe_mdb_in_7_ ),
    .Y(_03426_)
  );
  NAND2X1 _10695_ (
    .A(_03639_),
    .B(_03424_),
    .Y(_03427_)
  );
  AND2X1 _10696_ (
    .A(_03426_),
    .B(_03427_),
    .Y(_03428_)
  );
  NAND2X1 _10697_ (
    .A(execution_unit_0.inst_dext_7_ ),
    .B(_03877_),
    .Y(_03429_)
  );
  OAI21X1 _10698_ (
    .A(_03877_),
    .B(_03428_),
    .C(_03429_),
    .Y(_03354_)
  );
  NAND2X1 _10699_ (
    .A(execution_unit_0.inst_dext_8_ ),
    .B(_03877_),
    .Y(_03430_)
  );
  NAND3X1 _10700_ (
    .A(_03638_),
    .B(_03639_),
    .C(_03424_),
    .Y(_03431_)
  );
  XNOR2X1 _10701_ (
    .A(_03638_),
    .B(_03427_),
    .Y(_03432_)
  );
  OAI21X1 _10702_ (
    .A(_03877_),
    .B(_03432_),
    .C(_03430_),
    .Y(_03355_)
  );
  OAI21X1 _10703_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(_03427_),
    .C(dbg_0.fe_mdb_in_9_ ),
    .Y(_03433_)
  );
  OR2X1 _10704_ (
    .A(dbg_0.fe_mdb_in_9_ ),
    .B(_03431_),
    .Y(_03434_)
  );
  AND2X1 _10705_ (
    .A(_03433_),
    .B(_03434_),
    .Y(_03435_)
  );
  NAND2X1 _10706_ (
    .A(execution_unit_0.inst_dext_9_ ),
    .B(_03877_),
    .Y(_03436_)
  );
  OAI21X1 _10707_ (
    .A(_03877_),
    .B(_03435_),
    .C(_03436_),
    .Y(_03356_)
  );
  NAND2X1 _10708_ (
    .A(execution_unit_0.inst_dext_10_ ),
    .B(_03877_),
    .Y(_03437_)
  );
  NOR2X1 _10709_ (
    .A(dbg_0.fe_mdb_in_10_ ),
    .B(_03434_),
    .Y(_03438_)
  );
  XOR2X1 _10710_ (
    .A(dbg_0.fe_mdb_in_10_ ),
    .B(_03434_),
    .Y(_03439_)
  );
  OAI21X1 _10711_ (
    .A(_03877_),
    .B(_03439_),
    .C(_03437_),
    .Y(_03342_)
  );
  XNOR2X1 _10712_ (
    .A(dbg_0.fe_mdb_in_11_ ),
    .B(_03438_),
    .Y(_03440_)
  );
  NAND2X1 _10713_ (
    .A(execution_unit_0.inst_dext_11_ ),
    .B(_03877_),
    .Y(_03441_)
  );
  OAI21X1 _10714_ (
    .A(_03877_),
    .B(_03440_),
    .C(_03441_),
    .Y(_03343_)
  );
  NAND2X1 _10715_ (
    .A(execution_unit_0.inst_dext_12_ ),
    .B(_03877_),
    .Y(_03442_)
  );
  NOR2X1 _10716_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(dbg_0.fe_mdb_in_6_ ),
    .Y(_03443_)
  );
  NAND3X1 _10717_ (
    .A(_03752_),
    .B(_04073_),
    .C(_03443_),
    .Y(_03444_)
  );
  NOR2X1 _10718_ (
    .A(_03420_),
    .B(_03444_),
    .Y(_03445_)
  );
  OAI21X1 _10719_ (
    .A(_03420_),
    .B(_03444_),
    .C(dbg_0.fe_mdb_in_12_ ),
    .Y(_03446_)
  );
  NAND2X1 _10720_ (
    .A(_03673_),
    .B(_03445_),
    .Y(_03447_)
  );
  AND2X1 _10721_ (
    .A(_03446_),
    .B(_03447_),
    .Y(_03448_)
  );
  OAI21X1 _10722_ (
    .A(_03877_),
    .B(_03448_),
    .C(_03442_),
    .Y(_03344_)
  );
  OR2X1 _10723_ (
    .A(dbg_0.fe_mdb_in_13_ ),
    .B(_03447_),
    .Y(_03449_)
  );
  XNOR2X1 _10724_ (
    .A(_03640_),
    .B(_03447_),
    .Y(_03450_)
  );
  NAND2X1 _10725_ (
    .A(execution_unit_0.inst_dext_13_ ),
    .B(_03877_),
    .Y(_03451_)
  );
  OAI21X1 _10726_ (
    .A(_03877_),
    .B(_03450_),
    .C(_03451_),
    .Y(_03345_)
  );
  NAND2X1 _10727_ (
    .A(execution_unit_0.inst_dext_14_ ),
    .B(_03877_),
    .Y(_03452_)
  );
  NOR2X1 _10728_ (
    .A(dbg_0.fe_mdb_in_14_ ),
    .B(_03449_),
    .Y(_03453_)
  );
  XNOR2X1 _10729_ (
    .A(_03641_),
    .B(_03449_),
    .Y(_03454_)
  );
  OAI21X1 _10730_ (
    .A(_03877_),
    .B(_03454_),
    .C(_03452_),
    .Y(_03346_)
  );
  XNOR2X1 _10731_ (
    .A(dbg_0.fe_mdb_in_15_ ),
    .B(_03453_),
    .Y(_03455_)
  );
  NAND2X1 _10732_ (
    .A(execution_unit_0.inst_dext_15_ ),
    .B(_03877_),
    .Y(_03456_)
  );
  OAI21X1 _10733_ (
    .A(_03877_),
    .B(_03455_),
    .C(_03456_),
    .Y(_03347_)
  );
  NOR2X1 _10734_ (
    .A(_04037_),
    .B(_04106_),
    .Y(_03457_)
  );
  NAND2X1 _10735_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(_03457_),
    .Y(_03458_)
  );
  OAI21X1 _10736_ (
    .A(execution_unit_0.inst_sext_0_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03459_)
  );
  INVX1 _10737_ (
    .A(_03459_),
    .Y(_03460_)
  );
  OAI21X1 _10738_ (
    .A(dbg_0.fe_mdb_in_0_ ),
    .B(_03816_),
    .C(_03460_),
    .Y(_03461_)
  );
  OAI21X1 _10739_ (
    .A(_04108_),
    .B(_03461_),
    .C(_03458_),
    .Y(_03362_)
  );
  OAI21X1 _10740_ (
    .A(execution_unit_0.inst_sext_1_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03462_)
  );
  AOI21X1 _10741_ (
    .A(_03815_),
    .B(_03409_),
    .C(_03462_),
    .Y(_03463_)
  );
  AOI21X1 _10742_ (
    .A(dbg_0.fe_mdb_in_0_ ),
    .B(_04123_),
    .C(_03463_),
    .Y(_03464_)
  );
  NAND2X1 _10743_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_03457_),
    .Y(_03465_)
  );
  OAI21X1 _10744_ (
    .A(_04108_),
    .B(_03464_),
    .C(_03465_),
    .Y(_03369_)
  );
  NOR2X1 _10745_ (
    .A(_03761_),
    .B(_04104_),
    .Y(_03466_)
  );
  NOR2X1 _10746_ (
    .A(_03749_),
    .B(_03782_),
    .Y(_03467_)
  );
  NOR2X1 _10747_ (
    .A(_03466_),
    .B(_03467_),
    .Y(_03468_)
  );
  OAI21X1 _10748_ (
    .A(execution_unit_0.inst_sext_2_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03469_)
  );
  AOI21X1 _10749_ (
    .A(_03815_),
    .B(_03412_),
    .C(_03469_),
    .Y(_03470_)
  );
  AOI21X1 _10750_ (
    .A(dbg_0.fe_mdb_in_1_ ),
    .B(_04123_),
    .C(_03470_),
    .Y(_03471_)
  );
  MUX2X1 _10751_ (
    .A(_03468_),
    .B(_03471_),
    .S(_04108_),
    .Y(_03370_)
  );
  OAI21X1 _10752_ (
    .A(execution_unit_0.inst_sext_3_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03472_)
  );
  AOI21X1 _10753_ (
    .A(_03815_),
    .B(_03415_),
    .C(_03472_),
    .Y(_03473_)
  );
  AOI21X1 _10754_ (
    .A(dbg_0.fe_mdb_in_2_ ),
    .B(_04123_),
    .C(_03473_),
    .Y(_03474_)
  );
  MUX2X1 _10755_ (
    .A(_03749_),
    .B(_03474_),
    .S(_04108_),
    .Y(_03371_)
  );
  OAI21X1 _10756_ (
    .A(execution_unit_0.inst_sext_4_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03475_)
  );
  AOI21X1 _10757_ (
    .A(_03815_),
    .B(_03418_),
    .C(_03475_),
    .Y(_03476_)
  );
  AOI21X1 _10758_ (
    .A(dbg_0.fe_mdb_in_3_ ),
    .B(_04123_),
    .C(_03476_),
    .Y(_03477_)
  );
  NAND2X1 _10759_ (
    .A(_04108_),
    .B(_03467_),
    .Y(_03478_)
  );
  OAI21X1 _10760_ (
    .A(_04108_),
    .B(_03477_),
    .C(_03478_),
    .Y(_03372_)
  );
  OAI21X1 _10761_ (
    .A(execution_unit_0.inst_sext_5_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03479_)
  );
  AOI21X1 _10762_ (
    .A(_03815_),
    .B(_03421_),
    .C(_03479_),
    .Y(_03480_)
  );
  AOI21X1 _10763_ (
    .A(dbg_0.fe_mdb_in_4_ ),
    .B(_04123_),
    .C(_03480_),
    .Y(_03481_)
  );
  OAI21X1 _10764_ (
    .A(_04108_),
    .B(_03481_),
    .C(_03478_),
    .Y(_03373_)
  );
  OAI21X1 _10765_ (
    .A(execution_unit_0.inst_sext_6_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03482_)
  );
  AOI21X1 _10766_ (
    .A(_03815_),
    .B(_03425_),
    .C(_03482_),
    .Y(_03483_)
  );
  AOI21X1 _10767_ (
    .A(dbg_0.fe_mdb_in_5_ ),
    .B(_04123_),
    .C(_03483_),
    .Y(_03484_)
  );
  OAI21X1 _10768_ (
    .A(_04108_),
    .B(_03484_),
    .C(_03478_),
    .Y(_03374_)
  );
  OAI21X1 _10769_ (
    .A(execution_unit_0.inst_sext_7_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03485_)
  );
  AOI21X1 _10770_ (
    .A(_03815_),
    .B(_03428_),
    .C(_03485_),
    .Y(_03486_)
  );
  AOI21X1 _10771_ (
    .A(dbg_0.fe_mdb_in_6_ ),
    .B(_04123_),
    .C(_03486_),
    .Y(_03487_)
  );
  OAI21X1 _10772_ (
    .A(_04108_),
    .B(_03487_),
    .C(_03478_),
    .Y(_03375_)
  );
  OAI21X1 _10773_ (
    .A(execution_unit_0.inst_sext_8_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03488_)
  );
  AOI21X1 _10774_ (
    .A(_03815_),
    .B(_03432_),
    .C(_03488_),
    .Y(_03489_)
  );
  AOI21X1 _10775_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(_04123_),
    .C(_03489_),
    .Y(_03490_)
  );
  OAI21X1 _10776_ (
    .A(_04108_),
    .B(_03490_),
    .C(_03478_),
    .Y(_03376_)
  );
  OAI21X1 _10777_ (
    .A(execution_unit_0.inst_sext_9_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03491_)
  );
  AOI21X1 _10778_ (
    .A(_03815_),
    .B(_03435_),
    .C(_03491_),
    .Y(_03492_)
  );
  AOI21X1 _10779_ (
    .A(dbg_0.fe_mdb_in_8_ ),
    .B(_04123_),
    .C(_03492_),
    .Y(_03493_)
  );
  OAI21X1 _10780_ (
    .A(_04108_),
    .B(_03493_),
    .C(_03478_),
    .Y(_03377_)
  );
  OAI21X1 _10781_ (
    .A(execution_unit_0.inst_sext_10_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03494_)
  );
  AOI21X1 _10782_ (
    .A(_03815_),
    .B(_03439_),
    .C(_03494_),
    .Y(_03495_)
  );
  NOR2X1 _10783_ (
    .A(_03637_),
    .B(_04124_),
    .Y(_03496_)
  );
  NOR2X1 _10784_ (
    .A(_03495_),
    .B(_03496_),
    .Y(_03497_)
  );
  OAI21X1 _10785_ (
    .A(_04108_),
    .B(_03497_),
    .C(_03478_),
    .Y(_03363_)
  );
  OAI21X1 _10786_ (
    .A(execution_unit_0.inst_sext_11_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03498_)
  );
  AOI21X1 _10787_ (
    .A(_03815_),
    .B(_03440_),
    .C(_03498_),
    .Y(_03499_)
  );
  NOR2X1 _10788_ (
    .A(_03496_),
    .B(_03499_),
    .Y(_03500_)
  );
  OAI21X1 _10789_ (
    .A(_04108_),
    .B(_03500_),
    .C(_03478_),
    .Y(_03364_)
  );
  OAI21X1 _10790_ (
    .A(execution_unit_0.inst_sext_12_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03501_)
  );
  AOI21X1 _10791_ (
    .A(_03815_),
    .B(_03448_),
    .C(_03501_),
    .Y(_03502_)
  );
  NOR2X1 _10792_ (
    .A(_03496_),
    .B(_03502_),
    .Y(_03503_)
  );
  OAI21X1 _10793_ (
    .A(_04108_),
    .B(_03503_),
    .C(_03478_),
    .Y(_03365_)
  );
  OAI21X1 _10794_ (
    .A(execution_unit_0.inst_sext_13_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03504_)
  );
  AOI21X1 _10795_ (
    .A(_03815_),
    .B(_03450_),
    .C(_03504_),
    .Y(_03505_)
  );
  NOR2X1 _10796_ (
    .A(_03496_),
    .B(_03505_),
    .Y(_03506_)
  );
  OAI21X1 _10797_ (
    .A(_04108_),
    .B(_03506_),
    .C(_03478_),
    .Y(_03366_)
  );
  OAI21X1 _10798_ (
    .A(execution_unit_0.inst_sext_14_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03507_)
  );
  AOI21X1 _10799_ (
    .A(_03815_),
    .B(_03454_),
    .C(_03507_),
    .Y(_03508_)
  );
  NOR2X1 _10800_ (
    .A(_03496_),
    .B(_03508_),
    .Y(_03509_)
  );
  OAI21X1 _10801_ (
    .A(_04108_),
    .B(_03509_),
    .C(_03478_),
    .Y(_03367_)
  );
  OAI21X1 _10802_ (
    .A(execution_unit_0.inst_sext_15_ ),
    .B(_03815_),
    .C(_04124_),
    .Y(_03510_)
  );
  AOI21X1 _10803_ (
    .A(_03815_),
    .B(_03455_),
    .C(_03510_),
    .Y(_03511_)
  );
  NOR2X1 _10804_ (
    .A(_03496_),
    .B(_03511_),
    .Y(_03512_)
  );
  OAI21X1 _10805_ (
    .A(_04108_),
    .B(_03512_),
    .C(_03478_),
    .Y(_03368_)
  );
  NAND2X1 _10806_ (
    .A(_03633_),
    .B(_03717_),
    .Y(_03513_)
  );
  OR2X1 _10807_ (
    .A(irq_11_),
    .B(_03513_),
    .Y(_03514_)
  );
  NAND2X1 _10808_ (
    .A(irq_9_),
    .B(_03719_),
    .Y(_03515_)
  );
  OAI22X1 _10809_ (
    .A(1'h0),
    .B(_03717_),
    .C(_03514_),
    .D(_03515_),
    .Y(_03516_)
  );
  AOI21X1 _10810_ (
    .A(irq_12_),
    .B(_03628_),
    .C(1'h0),
    .Y(_03517_)
  );
  OAI21X1 _10811_ (
    .A(_03719_),
    .B(_03514_),
    .C(_03517_),
    .Y(_03518_)
  );
  AOI21X1 _10812_ (
    .A(_03719_),
    .B(_03720_),
    .C(_03513_),
    .Y(_03519_)
  );
  NOR2X1 _10813_ (
    .A(_03516_),
    .B(_03519_),
    .Y(_03520_)
  );
  NAND2X1 _10814_ (
    .A(irq_8_),
    .B(_03520_),
    .Y(_03521_)
  );
  NOR2X1 _10815_ (
    .A(_03518_),
    .B(_03521_),
    .Y(_03522_)
  );
  OR2X1 _10816_ (
    .A(_03516_),
    .B(_03522_),
    .Y(_03523_)
  );
  INVX1 _10817_ (
    .A(_03523_),
    .Y(_03524_)
  );
  AOI21X1 _10818_ (
    .A(irq_8_),
    .B(_03520_),
    .C(_03518_),
    .Y(_03525_)
  );
  NAND3X1 _10819_ (
    .A(irq_6_),
    .B(_03629_),
    .C(_03520_),
    .Y(_03526_)
  );
  AND2X1 _10820_ (
    .A(_03525_),
    .B(_03526_),
    .Y(_03527_)
  );
  INVX1 _10821_ (
    .A(_03527_),
    .Y(_03528_)
  );
  NOR2X1 _10822_ (
    .A(_03519_),
    .B(_03528_),
    .Y(_03529_)
  );
  NAND2X1 _10823_ (
    .A(irq_4_),
    .B(_03529_),
    .Y(_03530_)
  );
  NAND2X1 _10824_ (
    .A(irq_5_),
    .B(_03520_),
    .Y(_03531_)
  );
  NOR2X1 _10825_ (
    .A(_03522_),
    .B(_03531_),
    .Y(_03532_)
  );
  NAND2X1 _10826_ (
    .A(_03527_),
    .B(_03532_),
    .Y(_03533_)
  );
  NOR2X1 _10827_ (
    .A(_03523_),
    .B(_03530_),
    .Y(_03534_)
  );
  AND2X1 _10828_ (
    .A(_03520_),
    .B(_03525_),
    .Y(_03535_)
  );
  OAI21X1 _10829_ (
    .A(irq_6_),
    .B(irq_7_),
    .C(_03535_),
    .Y(_03536_)
  );
  NAND2X1 _10830_ (
    .A(_03533_),
    .B(_03536_),
    .Y(_03537_)
  );
  NAND3X1 _10831_ (
    .A(_03533_),
    .B(_03534_),
    .C(_03536_),
    .Y(_03538_)
  );
  NAND3X1 _10832_ (
    .A(_03527_),
    .B(_03532_),
    .C(_03536_),
    .Y(_03539_)
  );
  NAND3X1 _10833_ (
    .A(_03524_),
    .B(_03538_),
    .C(_03539_),
    .Y(_03540_)
  );
  NOR2X1 _10834_ (
    .A(_03534_),
    .B(_03537_),
    .Y(_03541_)
  );
  NAND2X1 _10835_ (
    .A(_03529_),
    .B(_03541_),
    .Y(_03542_)
  );
  NOR2X1 _10836_ (
    .A(_03540_),
    .B(_03542_),
    .Y(_03543_)
  );
  NAND3X1 _10837_ (
    .A(irq_2_),
    .B(_03630_),
    .C(_03543_),
    .Y(_03544_)
  );
  NAND3X1 _10838_ (
    .A(_03527_),
    .B(_03538_),
    .C(_03544_),
    .Y(_03545_)
  );
  NOR2X1 _10839_ (
    .A(_03734_),
    .B(_03545_),
    .Y(_03546_)
  );
  NAND2X1 _10840_ (
    .A(irq_3_),
    .B(_03543_),
    .Y(_03547_)
  );
  NOR2X1 _10841_ (
    .A(_03519_),
    .B(_03522_),
    .Y(_03548_)
  );
  NAND3X1 _10842_ (
    .A(_03544_),
    .B(_03547_),
    .C(_03548_),
    .Y(_03549_)
  );
  NOR2X1 _10843_ (
    .A(_03540_),
    .B(_03549_),
    .Y(_03550_)
  );
  NAND3X1 _10844_ (
    .A(_03541_),
    .B(_03544_),
    .C(_03547_),
    .Y(_03551_)
  );
  NOR2X1 _10845_ (
    .A(_03545_),
    .B(_03551_),
    .Y(_03552_)
  );
  AND2X1 _10846_ (
    .A(_03631_),
    .B(_03550_),
    .Y(_03553_)
  );
  NAND3X1 _10847_ (
    .A(irq_0_),
    .B(_03552_),
    .C(_03553_),
    .Y(_03554_)
  );
  NAND3X1 _10848_ (
    .A(irq_1_),
    .B(_03550_),
    .C(_03552_),
    .Y(_03555_)
  );
  NAND2X1 _10849_ (
    .A(_03546_),
    .B(_03554_),
    .Y(_03556_)
  );
  OAI21X1 _10850_ (
    .A(_03657_),
    .B(_03733_),
    .C(_03556_),
    .Y(_03394_)
  );
  NAND3X1 _10851_ (
    .A(_03733_),
    .B(_03554_),
    .C(_03555_),
    .Y(_03557_)
  );
  OAI22X1 _10852_ (
    .A(_03659_),
    .B(_03733_),
    .C(_03540_),
    .D(_03557_),
    .Y(_03395_)
  );
  OAI22X1 _10853_ (
    .A(_03661_),
    .B(_03733_),
    .C(_03549_),
    .D(_03557_),
    .Y(_03396_)
  );
  OAI21X1 _10854_ (
    .A(_03716_),
    .B(_03732_),
    .C(frontend_0.irq_addr_4_ ),
    .Y(_03558_)
  );
  OAI21X1 _10855_ (
    .A(_03551_),
    .B(_03557_),
    .C(_03558_),
    .Y(_03397_)
  );
  OR2X1 _10856_ (
    .A(frontend_0.irq_addr_5_ ),
    .B(_03733_),
    .Y(_03398_)
  );
  OAI21X1 _10857_ (
    .A(_03716_),
    .B(_03732_),
    .C(_03666_),
    .Y(_03399_)
  );
  NOR2X1 _10858_ (
    .A(_03696_),
    .B(exec_done),
    .Y(_03357_)
  );
  OAI21X1 _10859_ (
    .A(_03404_),
    .B(_03400_),
    .C(_03729_),
    .Y(_03559_)
  );
  NOR2X1 _10860_ (
    .A(_03841_),
    .B(_03559_),
    .Y(_03560_)
  );
  NAND2X1 _10861_ (
    .A(_04138_),
    .B(_03560_),
    .Y(_03561_)
  );
  INVX1 _10862_ (
    .A(_03561_),
    .Y(_03307_)
  );
  AND2X1 _10863_ (
    .A(frontend_0.irq_addr_5_ ),
    .B(frontend_0.irq_addr_6_ ),
    .Y(_03562_)
  );
  NAND2X1 _10864_ (
    .A(frontend_0.irq_addr_5_ ),
    .B(frontend_0.irq_addr_6_ ),
    .Y(_03563_)
  );
  NOR2X1 _10865_ (
    .A(_03657_),
    .B(frontend_0.irq_addr_2_ ),
    .Y(_03564_)
  );
  NAND2X1 _10866_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(_03659_),
    .Y(_03565_)
  );
  AND2X1 _10867_ (
    .A(frontend_0.irq_addr_3_ ),
    .B(frontend_0.irq_addr_4_ ),
    .Y(_03566_)
  );
  NAND2X1 _10868_ (
    .A(_03564_),
    .B(_03566_),
    .Y(_03567_)
  );
  NAND2X1 _10869_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(frontend_0.irq_addr_2_ ),
    .Y(_03568_)
  );
  INVX1 _10870_ (
    .A(_03568_),
    .Y(_03569_)
  );
  NAND2X1 _10871_ (
    .A(_03661_),
    .B(frontend_0.irq_addr_4_ ),
    .Y(_03570_)
  );
  OAI21X1 _10872_ (
    .A(_03568_),
    .B(_03570_),
    .C(_03567_),
    .Y(_03571_)
  );
  NAND2X1 _10873_ (
    .A(_03562_),
    .B(_03571_),
    .Y(_03572_)
  );
  NAND3X1 _10874_ (
    .A(_03562_),
    .B(_03565_),
    .C(_03566_),
    .Y(_03573_)
  );
  NOR2X1 _10875_ (
    .A(_03563_),
    .B(_03570_),
    .Y(_03574_)
  );
  OR2X1 _10876_ (
    .A(_03563_),
    .B(_03570_),
    .Y(_03575_)
  );
  NOR2X1 _10877_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(frontend_0.irq_addr_2_ ),
    .Y(_03576_)
  );
  INVX1 _10878_ (
    .A(_03576_),
    .Y(_03577_)
  );
  NOR2X1 _10879_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(_03659_),
    .Y(_03578_)
  );
  NAND2X1 _10880_ (
    .A(_03657_),
    .B(frontend_0.irq_addr_2_ ),
    .Y(_03579_)
  );
  OAI21X1 _10881_ (
    .A(_03564_),
    .B(_03578_),
    .C(_03574_),
    .Y(_03580_)
  );
  NAND3X1 _10882_ (
    .A(_03572_),
    .B(_03573_),
    .C(_03580_),
    .Y(_03581_)
  );
  OR2X1 _10883_ (
    .A(_03570_),
    .B(_03577_),
    .Y(_03582_)
  );
  NOR2X1 _10884_ (
    .A(_03661_),
    .B(frontend_0.irq_addr_4_ ),
    .Y(_03583_)
  );
  OAI21X1 _10885_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(frontend_0.irq_addr_2_ ),
    .C(_03583_),
    .Y(_03584_)
  );
  AOI21X1 _10886_ (
    .A(_03582_),
    .B(_03584_),
    .C(_03563_),
    .Y(_03585_)
  );
  OR2X1 _10887_ (
    .A(_03581_),
    .B(_03585_),
    .Y(_03586_)
  );
  NOR2X1 _10888_ (
    .A(frontend_0.irq_addr_3_ ),
    .B(frontend_0.irq_addr_4_ ),
    .Y(_03587_)
  );
  AOI22X1 _10889_ (
    .A(_03576_),
    .B(_03583_),
    .C(_03587_),
    .D(_03569_),
    .Y(_03588_)
  );
  NOR2X1 _10890_ (
    .A(_03666_),
    .B(_03921_),
    .Y(_03589_)
  );
  OR2X1 _10891_ (
    .A(_03666_),
    .B(_03921_),
    .Y(_03590_)
  );
  OAI21X1 _10892_ (
    .A(_03564_),
    .B(_03578_),
    .C(_03587_),
    .Y(_03591_)
  );
  AND2X1 _10893_ (
    .A(_03589_),
    .B(_03591_),
    .Y(_03592_)
  );
  OAI21X1 _10894_ (
    .A(_03563_),
    .B(_03588_),
    .C(_03592_),
    .Y(_03593_)
  );
  NOR2X1 _10895_ (
    .A(_03586_),
    .B(_03593_),
    .Y(_00083_)
  );
  OR2X1 _10896_ (
    .A(_03586_),
    .B(_03590_),
    .Y(_03594_)
  );
  INVX1 _10897_ (
    .A(_03594_),
    .Y(_03595_)
  );
  NAND2X1 _10898_ (
    .A(_03588_),
    .B(_03595_),
    .Y(_03596_)
  );
  AOI21X1 _10899_ (
    .A(_03657_),
    .B(_03587_),
    .C(_03596_),
    .Y(_00088_)
  );
  NAND2X1 _10900_ (
    .A(_03562_),
    .B(_03587_),
    .Y(_03597_)
  );
  NOR2X1 _10901_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03597_),
    .Y(_03598_)
  );
  NOR2X1 _10902_ (
    .A(_03596_),
    .B(_03598_),
    .Y(_00089_)
  );
  AOI22X1 _10903_ (
    .A(_03576_),
    .B(_03583_),
    .C(_03587_),
    .D(_03578_),
    .Y(_03599_)
  );
  OAI21X1 _10904_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03597_),
    .C(_03599_),
    .Y(_03600_)
  );
  NOR2X1 _10905_ (
    .A(_03594_),
    .B(_03600_),
    .Y(_00090_)
  );
  NOR2X1 _10906_ (
    .A(_03587_),
    .B(_03594_),
    .Y(_00091_)
  );
  NAND3X1 _10907_ (
    .A(_03582_),
    .B(_03589_),
    .C(_03597_),
    .Y(_03601_)
  );
  OR2X1 _10908_ (
    .A(_03581_),
    .B(_03601_),
    .Y(_03602_)
  );
  AOI21X1 _10909_ (
    .A(_03565_),
    .B(_03583_),
    .C(_03602_),
    .Y(_00092_)
  );
  OAI21X1 _10910_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03563_),
    .C(_03568_),
    .Y(_03603_)
  );
  AOI21X1 _10911_ (
    .A(_03583_),
    .B(_03603_),
    .C(_03602_),
    .Y(_00093_)
  );
  OAI21X1 _10912_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03563_),
    .C(_03579_),
    .Y(_03604_)
  );
  AOI21X1 _10913_ (
    .A(_03583_),
    .B(_03604_),
    .C(_03602_),
    .Y(_00094_)
  );
  NAND3X1 _10914_ (
    .A(frontend_0.irq_addr_4_ ),
    .B(_03573_),
    .C(_03589_),
    .Y(_03605_)
  );
  INVX1 _10915_ (
    .A(_03605_),
    .Y(_03606_)
  );
  NOR2X1 _10916_ (
    .A(_03571_),
    .B(_03605_),
    .Y(_03607_)
  );
  AND2X1 _10917_ (
    .A(_03580_),
    .B(_03607_),
    .Y(_00095_)
  );
  OAI21X1 _10918_ (
    .A(frontend_0.irq_addr_1_ ),
    .B(_03575_),
    .C(_03607_),
    .Y(_03608_)
  );
  INVX1 _10919_ (
    .A(_03608_),
    .Y(_00096_)
  );
  OAI21X1 _10920_ (
    .A(frontend_0.irq_addr_2_ ),
    .B(_03575_),
    .C(_03606_),
    .Y(_03609_)
  );
  AOI21X1 _10921_ (
    .A(_03562_),
    .B(_03571_),
    .C(_03609_),
    .Y(_00084_)
  );
  OAI21X1 _10922_ (
    .A(_03570_),
    .B(_03579_),
    .C(_03567_),
    .Y(_03610_)
  );
  AOI21X1 _10923_ (
    .A(_03562_),
    .B(_03610_),
    .C(_03609_),
    .Y(_00085_)
  );
  NAND2X1 _10924_ (
    .A(_03566_),
    .B(_03589_),
    .Y(_03611_)
  );
  NOR2X1 _10925_ (
    .A(_03577_),
    .B(_03611_),
    .Y(_00086_)
  );
  NOR2X1 _10926_ (
    .A(_03567_),
    .B(_03590_),
    .Y(_00087_)
  );
  OR2X1 _10927_ (
    .A(frontend_0.pmem_busy ),
    .B(_03849_),
    .Y(_03612_)
  );
  AOI21X1 _10928_ (
    .A(cpu_halt_st),
    .B(_03728_),
    .C(_03612_),
    .Y(_03613_)
  );
  OAI21X1 _10929_ (
    .A(_03830_),
    .B(_03887_),
    .C(_03613_),
    .Y(fe_mb_en)
  );
  OR2X1 _10930_ (
    .A(_03681_),
    .B(frontend_0.inst_jmp_bin_2_ ),
    .Y(_03614_)
  );
  NAND2X1 _10931_ (
    .A(_03694_),
    .B(_03695_),
    .Y(_03615_)
  );
  NOR2X1 _10932_ (
    .A(_03614_),
    .B(_03615_),
    .Y(execution_unit_0.alu_0.inst_jmp_0_ )
  );
  NAND2X1 _10933_ (
    .A(frontend_0.inst_jmp_bin_0_ ),
    .B(_03695_),
    .Y(_03616_)
  );
  NOR2X1 _10934_ (
    .A(_03614_),
    .B(_03616_),
    .Y(execution_unit_0.alu_0.inst_jmp_1_ )
  );
  NAND2X1 _10935_ (
    .A(_03694_),
    .B(frontend_0.inst_jmp_bin_1_ ),
    .Y(_03617_)
  );
  NOR2X1 _10936_ (
    .A(_03614_),
    .B(_03617_),
    .Y(execution_unit_0.alu_0.inst_jmp_2_ )
  );
  NAND2X1 _10937_ (
    .A(frontend_0.inst_jmp_bin_0_ ),
    .B(frontend_0.inst_jmp_bin_1_ ),
    .Y(_03618_)
  );
  NOR2X1 _10938_ (
    .A(_03614_),
    .B(_03618_),
    .Y(execution_unit_0.alu_0.inst_jmp_3_ )
  );
  NAND2X1 _10939_ (
    .A(execution_unit_0.inst_type_1_ ),
    .B(frontend_0.inst_jmp_bin_2_ ),
    .Y(_03619_)
  );
  NOR2X1 _10940_ (
    .A(_03615_),
    .B(_03619_),
    .Y(execution_unit_0.alu_0.inst_jmp_4_ )
  );
  NOR2X1 _10941_ (
    .A(_03616_),
    .B(_03619_),
    .Y(execution_unit_0.alu_0.inst_jmp_5_ )
  );
  NOR2X1 _10942_ (
    .A(_03617_),
    .B(_03619_),
    .Y(execution_unit_0.alu_0.inst_jmp_6_ )
  );
  NAND2X1 _10943_ (
    .A(execution_unit_0.inst_type_0_ ),
    .B(_03804_),
    .Y(_03620_)
  );
  OAI21X1 _10944_ (
    .A(_03703_),
    .B(_03704_),
    .C(frontend_0.exec_src_wr ),
    .Y(_03621_)
  );
  OAI21X1 _10945_ (
    .A(_03711_),
    .B(_03621_),
    .C(_03620_),
    .Y(_03311_)
  );
  OAI21X1 _10946_ (
    .A(_03703_),
    .B(_03795_),
    .C(_03707_),
    .Y(_03309_)
  );
  NOR2X1 _10947_ (
    .A(dbg_0.fe_mdb_in_7_ ),
    .B(_04085_),
    .Y(_03622_)
  );
  AOI21X1 _10948_ (
    .A(_03773_),
    .B(_03622_),
    .C(_04058_),
    .Y(_03623_)
  );
  OAI21X1 _10949_ (
    .A(_04037_),
    .B(_03623_),
    .C(_03700_),
    .Y(_03310_)
  );
  DFFSR _10950_ (
    .CLK(dco_clk),
    .D(_03402_),
    .Q(frontend_0.i_state_0_ ),
    .R(1'h1),
    .S(_03405_)
  );
  DFFSR _10951_ (
    .CLK(dco_clk),
    .D(_03400_),
    .Q(frontend_0.i_state_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10952_ (
    .CLK(dco_clk),
    .D(_03403_),
    .Q(frontend_0.i_state_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10953_ (
    .CLK(dco_clk),
    .D(frontend_0.i_state_0_ ),
    .Q(frontend_0.i_state_3_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10954_ (
    .CLK(dco_clk),
    .D(_03404_),
    .Q(frontend_0.i_state_4_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10955_ (
    .CLK(dco_clk),
    .D(_03401_),
    .Q(frontend_0.i_state_5_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10956_ (
    .CLK(dco_clk),
    .D(_03316_),
    .Q(execution_unit_0.alu_0.inst_alu_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10957_ (
    .CLK(dco_clk),
    .D(_03319_),
    .Q(execution_unit_0.alu_0.inst_alu_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10958_ (
    .CLK(dco_clk),
    .D(_03320_),
    .Q(execution_unit_0.alu_0.inst_alu_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10959_ (
    .CLK(dco_clk),
    .D(_03321_),
    .Q(execution_unit_0.alu_0.inst_alu_3_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10960_ (
    .CLK(dco_clk),
    .D(_03322_),
    .Q(execution_unit_0.alu_0.inst_alu_4_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10961_ (
    .CLK(dco_clk),
    .D(_03323_),
    .Q(execution_unit_0.alu_0.inst_alu_5_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10962_ (
    .CLK(dco_clk),
    .D(_03324_),
    .Q(execution_unit_0.alu_0.inst_alu_6_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10963_ (
    .CLK(dco_clk),
    .D(_03325_),
    .Q(execution_unit_0.alu_0.inst_alu_7_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10964_ (
    .CLK(dco_clk),
    .D(_03326_),
    .Q(execution_unit_0.alu_0.inst_alu_8_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10965_ (
    .CLK(dco_clk),
    .D(_03327_),
    .Q(execution_unit_0.alu_0.inst_alu_9_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10966_ (
    .CLK(dco_clk),
    .D(_03317_),
    .Q(execution_unit_0.alu_0.inst_alu_10_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10967_ (
    .CLK(dco_clk),
    .D(_03318_),
    .Q(execution_unit_0.alu_0.UNUSED_inst_alu ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10968_ (
    .CLK(dco_clk),
    .D(frontend_0.e_state_nxt_0_ ),
    .Q(e_state_0_),
    .R(1'h1),
    .S(_03405_)
  );
  DFFSR _10969_ (
    .CLK(dco_clk),
    .D(frontend_0.e_state_nxt_1_ ),
    .Q(e_state_1_),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10970_ (
    .CLK(dco_clk),
    .D(frontend_0.e_state_nxt_2_ ),
    .Q(e_state_2_),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10971_ (
    .CLK(dco_clk),
    .D(frontend_0.e_state_nxt_3_ ),
    .Q(e_state_3_),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10972_ (
    .CLK(dco_clk),
    .D(_03308_),
    .Q(frontend_0.exec_dext_rdy ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10973_ (
    .CLK(dco_clk),
    .D(_03311_),
    .Q(frontend_0.exec_src_wr ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10974_ (
    .CLK(dco_clk),
    .D(_03309_),
    .Q(frontend_0.exec_dst_wr ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10975_ (
    .CLK(dco_clk),
    .D(_03310_),
    .Q(frontend_0.exec_jmp ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10976_ (
    .CLK(dco_clk),
    .D(_03389_),
    .Q(frontend_0.inst_sz_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10977_ (
    .CLK(dco_clk),
    .D(_03390_),
    .Q(frontend_0.inst_sz_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10978_ (
    .CLK(dco_clk),
    .D(_03336_),
    .Q(execution_unit_0.alu_0.inst_bw ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10979_ (
    .CLK(dco_clk),
    .D(_03312_),
    .Q(execution_unit_0.inst_ad_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10980_ (
    .CLK(dco_clk),
    .D(_03313_),
    .Q(execution_unit_0.UNUSED_inst_ad_idx ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10981_ (
    .CLK(dco_clk),
    .D(_03314_),
    .Q(execution_unit_0.UNUSED_inst_ad_symb ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10982_ (
    .CLK(dco_clk),
    .D(_03315_),
    .Q(execution_unit_0.inst_ad_6_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10983_ (
    .CLK(dco_clk),
    .D(_03328_),
    .Q(execution_unit_0.inst_as_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10984_ (
    .CLK(dco_clk),
    .D(_03329_),
    .Q(execution_unit_0.inst_as_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10985_ (
    .CLK(dco_clk),
    .D(_03330_),
    .Q(execution_unit_0.inst_as_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10986_ (
    .CLK(dco_clk),
    .D(_03331_),
    .Q(execution_unit_0.inst_as_3_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10987_ (
    .CLK(dco_clk),
    .D(_03332_),
    .Q(execution_unit_0.inst_as_4_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10988_ (
    .CLK(dco_clk),
    .D(_03333_),
    .Q(execution_unit_0.inst_as_5_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10989_ (
    .CLK(dco_clk),
    .D(_03334_),
    .Q(execution_unit_0.inst_as_6_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10990_ (
    .CLK(dco_clk),
    .D(_03335_),
    .Q(execution_unit_0.inst_as_7_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10991_ (
    .CLK(dco_clk),
    .D(_03385_),
    .Q(frontend_0.inst_src_bin_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10992_ (
    .CLK(dco_clk),
    .D(_03386_),
    .Q(frontend_0.inst_src_bin_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10993_ (
    .CLK(dco_clk),
    .D(_03387_),
    .Q(frontend_0.inst_src_bin_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10994_ (
    .CLK(dco_clk),
    .D(_03388_),
    .Q(frontend_0.inst_src_bin_3_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10995_ (
    .CLK(dco_clk),
    .D(_03337_),
    .Q(frontend_0.inst_dest_bin_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10996_ (
    .CLK(dco_clk),
    .D(_03338_),
    .Q(frontend_0.inst_dest_bin_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10997_ (
    .CLK(dco_clk),
    .D(_03339_),
    .Q(frontend_0.inst_dest_bin_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10998_ (
    .CLK(dco_clk),
    .D(_03340_),
    .Q(frontend_0.inst_dest_bin_3_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _10999_ (
    .CLK(dco_clk),
    .D(_03361_),
    .Q(execution_unit_0.inst_mov ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11000_ (
    .CLK(dco_clk),
    .D(_03358_),
    .Q(frontend_0.inst_jmp_bin_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11001_ (
    .CLK(dco_clk),
    .D(_03359_),
    .Q(frontend_0.inst_jmp_bin_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11002_ (
    .CLK(dco_clk),
    .D(_03360_),
    .Q(frontend_0.inst_jmp_bin_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11003_ (
    .CLK(dco_clk),
    .D(_03378_),
    .Q(execution_unit_0.alu_0.inst_so_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11004_ (
    .CLK(dco_clk),
    .D(_03379_),
    .Q(execution_unit_0.alu_0.inst_so_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11005_ (
    .CLK(dco_clk),
    .D(_03380_),
    .Q(execution_unit_0.alu_0.inst_so_3_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11006_ (
    .CLK(dco_clk),
    .D(_03381_),
    .Q(execution_unit_0.alu_0.UNUSED_inst_so_push ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11007_ (
    .CLK(dco_clk),
    .D(_03382_),
    .Q(execution_unit_0.alu_0.UNUSED_inst_so_call ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11008_ (
    .CLK(dco_clk),
    .D(_03383_),
    .Q(execution_unit_0.alu_0.UNUSED_inst_so_reti ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11009_ (
    .CLK(dco_clk),
    .D(_03384_),
    .Q(execution_unit_0.alu_0.inst_so_7_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11010_ (
    .CLK(dco_clk),
    .D(_03391_),
    .Q(execution_unit_0.inst_type_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11011_ (
    .CLK(dco_clk),
    .D(_03392_),
    .Q(execution_unit_0.inst_type_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11012_ (
    .CLK(dco_clk),
    .D(_03393_),
    .Q(execution_unit_0.inst_type_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11013_ (
    .CLK(dco_clk),
    .D(_03341_),
    .Q(execution_unit_0.inst_dext_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11014_ (
    .CLK(dco_clk),
    .D(_03348_),
    .Q(execution_unit_0.inst_dext_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11015_ (
    .CLK(dco_clk),
    .D(_03349_),
    .Q(execution_unit_0.inst_dext_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11016_ (
    .CLK(dco_clk),
    .D(_03350_),
    .Q(execution_unit_0.inst_dext_3_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11017_ (
    .CLK(dco_clk),
    .D(_03351_),
    .Q(execution_unit_0.inst_dext_4_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11018_ (
    .CLK(dco_clk),
    .D(_03352_),
    .Q(execution_unit_0.inst_dext_5_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11019_ (
    .CLK(dco_clk),
    .D(_03353_),
    .Q(execution_unit_0.inst_dext_6_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11020_ (
    .CLK(dco_clk),
    .D(_03354_),
    .Q(execution_unit_0.inst_dext_7_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11021_ (
    .CLK(dco_clk),
    .D(_03355_),
    .Q(execution_unit_0.inst_dext_8_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11022_ (
    .CLK(dco_clk),
    .D(_03356_),
    .Q(execution_unit_0.inst_dext_9_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11023_ (
    .CLK(dco_clk),
    .D(_03342_),
    .Q(execution_unit_0.inst_dext_10_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11024_ (
    .CLK(dco_clk),
    .D(_03343_),
    .Q(execution_unit_0.inst_dext_11_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11025_ (
    .CLK(dco_clk),
    .D(_03344_),
    .Q(execution_unit_0.inst_dext_12_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11026_ (
    .CLK(dco_clk),
    .D(_03345_),
    .Q(execution_unit_0.inst_dext_13_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11027_ (
    .CLK(dco_clk),
    .D(_03346_),
    .Q(execution_unit_0.inst_dext_14_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11028_ (
    .CLK(dco_clk),
    .D(_03347_),
    .Q(execution_unit_0.inst_dext_15_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11029_ (
    .CLK(dco_clk),
    .D(_03362_),
    .Q(execution_unit_0.inst_sext_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11030_ (
    .CLK(dco_clk),
    .D(_03369_),
    .Q(execution_unit_0.inst_sext_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11031_ (
    .CLK(dco_clk),
    .D(_03370_),
    .Q(execution_unit_0.inst_sext_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11032_ (
    .CLK(dco_clk),
    .D(_03371_),
    .Q(execution_unit_0.inst_sext_3_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11033_ (
    .CLK(dco_clk),
    .D(_03372_),
    .Q(execution_unit_0.inst_sext_4_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11034_ (
    .CLK(dco_clk),
    .D(_03373_),
    .Q(execution_unit_0.inst_sext_5_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11035_ (
    .CLK(dco_clk),
    .D(_03374_),
    .Q(execution_unit_0.inst_sext_6_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11036_ (
    .CLK(dco_clk),
    .D(_03375_),
    .Q(execution_unit_0.inst_sext_7_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11037_ (
    .CLK(dco_clk),
    .D(_03376_),
    .Q(execution_unit_0.inst_sext_8_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11038_ (
    .CLK(dco_clk),
    .D(_03377_),
    .Q(execution_unit_0.inst_sext_9_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11039_ (
    .CLK(dco_clk),
    .D(_03363_),
    .Q(execution_unit_0.inst_sext_10_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11040_ (
    .CLK(dco_clk),
    .D(_03364_),
    .Q(execution_unit_0.inst_sext_11_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11041_ (
    .CLK(dco_clk),
    .D(_03365_),
    .Q(execution_unit_0.inst_sext_12_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11042_ (
    .CLK(dco_clk),
    .D(_03366_),
    .Q(execution_unit_0.inst_sext_13_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11043_ (
    .CLK(dco_clk),
    .D(_03367_),
    .Q(execution_unit_0.inst_sext_14_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11044_ (
    .CLK(dco_clk),
    .D(_03368_),
    .Q(execution_unit_0.inst_sext_15_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11045_ (
    .CLK(dco_clk),
    .D(fe_pmem_wait),
    .Q(frontend_0.pmem_busy ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11046_ (
    .CLK(dco_clk),
    .D(UNUSED_fe_mab_0),
    .Q(dbg_0.UNUSED_pc_0_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11047_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_1_ ),
    .Q(dbg_0.UNUSED_pc_1_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11048_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_2_ ),
    .Q(dbg_0.UNUSED_pc_2_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11049_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_3_ ),
    .Q(dbg_0.UNUSED_pc_3_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11050_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_4_ ),
    .Q(dbg_0.UNUSED_pc_4_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11051_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_5_ ),
    .Q(dbg_0.UNUSED_pc_5_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11052_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_6_ ),
    .Q(dbg_0.UNUSED_pc_6_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11053_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_7_ ),
    .Q(dbg_0.UNUSED_pc_7_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11054_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_8_ ),
    .Q(dbg_0.UNUSED_pc_8_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11055_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_9_ ),
    .Q(dbg_0.UNUSED_pc_9_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11056_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_10_ ),
    .Q(dbg_0.UNUSED_pc_10_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11057_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_11_ ),
    .Q(dbg_0.UNUSED_pc_11_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11058_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_12_ ),
    .Q(dbg_0.UNUSED_pc_12_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11059_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_13_ ),
    .Q(dbg_0.UNUSED_pc_13_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11060_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_14_ ),
    .Q(dbg_0.UNUSED_pc_14_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11061_ (
    .CLK(dco_clk),
    .D(execution_unit_0.pc_nxt_15_ ),
    .Q(dbg_0.UNUSED_pc_15_ ),
    .R(_03405_),
    .S(1'h1)
  );
  DFFSR _11062_ (
    .CLK(dco_clk),
    .D(_03394_),
    .Q(frontend_0.irq_addr_1_ ),
    .R(1'h1),
    .S(_03405_)
  );
  DFFSR _11063_ (
    .CLK(dco_clk),
    .D(_03395_),
    .Q(frontend_0.irq_addr_2_ ),
    .R(1'h1),
    .S(_03405_)
  );
  DFFSR _11064_ (
    .CLK(dco_clk),
    .D(_03396_),
    .Q(frontend_0.irq_addr_3_ ),
    .R(1'h1),
    .S(_03405_)
  );
  DFFSR _11065_ (
    .CLK(dco_clk),
    .D(_03397_),
    .Q(frontend_0.irq_addr_4_ ),
    .R(1'h1),
    .S(_03405_)
  );
  DFFSR _11066_ (
    .CLK(dco_clk),
    .D(_03398_),
    .Q(frontend_0.irq_addr_5_ ),
    .R(1'h1),
    .S(_03405_)
  );
  DFFSR _11067_ (
    .CLK(dco_clk),
    .D(_03399_),
    .Q(frontend_0.irq_addr_6_ ),
    .R(1'h1),
    .S(_03405_)
  );
  DFFSR _11068_ (
    .CLK(dco_clk),
    .D(_03357_),
    .Q(execution_unit_0.inst_irq_rst ),
    .R(1'h1),
    .S(_03405_)
  );
  DFFSR _11069_ (
    .CLK(dco_clk),
    .D(_03307_),
    .Q(cpu_halt_st),
    .R(_03405_),
    .S(1'h1)
  );
  INVX1 _11070_ (
    .A(cpu_halt_st),
    .Y(_04166_)
  );
  INVX1 _11071_ (
    .A(pmem_dout_0_),
    .Y(_04167_)
  );
  INVX1 _11072_ (
    .A(pmem_dout_1_),
    .Y(_04168_)
  );
  INVX1 _11073_ (
    .A(pmem_dout_2_),
    .Y(_04169_)
  );
  INVX1 _11074_ (
    .A(pmem_dout_3_),
    .Y(_04170_)
  );
  INVX1 _11075_ (
    .A(pmem_dout_4_),
    .Y(_04171_)
  );
  INVX1 _11076_ (
    .A(pmem_dout_5_),
    .Y(_04172_)
  );
  INVX1 _11077_ (
    .A(pmem_dout_6_),
    .Y(_04173_)
  );
  INVX1 _11078_ (
    .A(pmem_dout_7_),
    .Y(_04174_)
  );
  INVX1 _11079_ (
    .A(pmem_dout_8_),
    .Y(_04175_)
  );
  INVX1 _11080_ (
    .A(pmem_dout_9_),
    .Y(_04176_)
  );
  INVX1 _11081_ (
    .A(pmem_dout_10_),
    .Y(_04177_)
  );
  INVX1 _11082_ (
    .A(pmem_dout_11_),
    .Y(_04178_)
  );
  INVX1 _11083_ (
    .A(pmem_dout_12_),
    .Y(_04179_)
  );
  INVX1 _11084_ (
    .A(pmem_dout_13_),
    .Y(_04180_)
  );
  INVX1 _11085_ (
    .A(pmem_dout_14_),
    .Y(_04181_)
  );
  INVX1 _11086_ (
    .A(pmem_dout_15_),
    .Y(_04182_)
  );
  INVX1 _11087_ (
    .A(dbg_0.UNUSED_eu_mb_wr_0_ ),
    .Y(_04183_)
  );
  INVX1 _11088_ (
    .A(dbg_0.dbg_mem_wr_0_ ),
    .Y(_04184_)
  );
  INVX1 _11089_ (
    .A(dbg_0.dbg_mem_addr_15_ ),
    .Y(_04185_)
  );
  INVX1 _11090_ (
    .A(dbg_0.dbg_mem_addr_14_ ),
    .Y(_04186_)
  );
  INVX1 _11091_ (
    .A(dbg_0.dbg_mem_addr_13_ ),
    .Y(_04187_)
  );
  INVX1 _11092_ (
    .A(dbg_0.dbg_mem_addr_12_ ),
    .Y(_04188_)
  );
  INVX1 _11093_ (
    .A(dbg_0.dbg_mem_addr_11_ ),
    .Y(_04189_)
  );
  INVX1 _11094_ (
    .A(dbg_0.dbg_mem_addr_10_ ),
    .Y(_04190_)
  );
  INVX1 _11095_ (
    .A(dbg_0.dbg_mem_addr_9_ ),
    .Y(_04191_)
  );
  INVX1 _11096_ (
    .A(dbg_0.dbg_mem_addr_8_ ),
    .Y(_04192_)
  );
  INVX1 _11097_ (
    .A(dbg_0.dbg_mem_addr_7_ ),
    .Y(_04193_)
  );
  INVX1 _11098_ (
    .A(dbg_0.dbg_mem_addr_6_ ),
    .Y(_04194_)
  );
  INVX1 _11099_ (
    .A(dbg_0.dbg_mem_addr_5_ ),
    .Y(_04195_)
  );
  INVX1 _11100_ (
    .A(dbg_0.dbg_mem_addr_4_ ),
    .Y(_04196_)
  );
  INVX1 _11101_ (
    .A(dbg_0.dbg_mem_addr_3_ ),
    .Y(_04197_)
  );
  INVX1 _11102_ (
    .A(dbg_0.dbg_mem_addr_2_ ),
    .Y(_04198_)
  );
  INVX1 _11103_ (
    .A(dbg_0.dbg_mem_addr_1_ ),
    .Y(_04199_)
  );
  INVX1 _11104_ (
    .A(dbg_0.UNUSED_eu_mb_en ),
    .Y(_04200_)
  );
  INVX1 _11105_ (
    .A(dbg_0.UNUSED_eu_mab_13_ ),
    .Y(_04201_)
  );
  INVX1 _11106_ (
    .A(dbg_0.UNUSED_eu_mab_12_ ),
    .Y(_04202_)
  );
  INVX1 _11107_ (
    .A(dbg_0.UNUSED_eu_mab_11_ ),
    .Y(_04203_)
  );
  INVX1 _11108_ (
    .A(dbg_0.UNUSED_eu_mab_10_ ),
    .Y(_04204_)
  );
  INVX1 _11109_ (
    .A(dbg_0.UNUSED_eu_mab_9_ ),
    .Y(_04205_)
  );
  INVX1 _11110_ (
    .A(dbg_0.UNUSED_eu_mab_8_ ),
    .Y(_04206_)
  );
  INVX1 _11111_ (
    .A(dbg_0.UNUSED_eu_mab_7_ ),
    .Y(_04207_)
  );
  INVX1 _11112_ (
    .A(dbg_0.UNUSED_eu_mab_6_ ),
    .Y(_04208_)
  );
  INVX1 _11113_ (
    .A(dbg_0.UNUSED_eu_mab_5_ ),
    .Y(_04209_)
  );
  INVX1 _11114_ (
    .A(dbg_0.UNUSED_eu_mab_4_ ),
    .Y(_04210_)
  );
  INVX1 _11115_ (
    .A(dbg_0.UNUSED_eu_mab_3_ ),
    .Y(_04211_)
  );
  INVX1 _11116_ (
    .A(dbg_0.UNUSED_eu_mab_2_ ),
    .Y(_04212_)
  );
  INVX1 _11117_ (
    .A(dbg_0.UNUSED_eu_mab_1_ ),
    .Y(_04213_)
  );
  INVX1 _11118_ (
    .A(dbg_0.UNUSED_eu_mb_wr_1_ ),
    .Y(_04214_)
  );
  INVX1 _11119_ (
    .A(dbg_0.dbg_mem_wr_1_ ),
    .Y(_04215_)
  );
  INVX1 _11120_ (
    .A(_00144_),
    .Y(_04216_)
  );
  INVX1 _11121_ (
    .A(eu_mdb_out_0_),
    .Y(_04217_)
  );
  INVX1 _11122_ (
    .A(_00151_),
    .Y(_04218_)
  );
  INVX1 _11123_ (
    .A(eu_mdb_out_1_),
    .Y(_04219_)
  );
  INVX1 _11124_ (
    .A(_00152_),
    .Y(_04220_)
  );
  INVX1 _11125_ (
    .A(eu_mdb_out_2_),
    .Y(_04221_)
  );
  INVX1 _11126_ (
    .A(_00153_),
    .Y(_04222_)
  );
  INVX1 _11127_ (
    .A(eu_mdb_out_3_),
    .Y(_04223_)
  );
  INVX1 _11128_ (
    .A(_00154_),
    .Y(_04224_)
  );
  INVX1 _11129_ (
    .A(eu_mdb_out_4_),
    .Y(_04225_)
  );
  INVX1 _11130_ (
    .A(_00155_),
    .Y(_04226_)
  );
  INVX1 _11131_ (
    .A(eu_mdb_out_5_),
    .Y(_04227_)
  );
  INVX1 _11132_ (
    .A(_00156_),
    .Y(_04228_)
  );
  INVX1 _11133_ (
    .A(eu_mdb_out_6_),
    .Y(_04229_)
  );
  INVX1 _11134_ (
    .A(_00157_),
    .Y(_04230_)
  );
  INVX1 _11135_ (
    .A(eu_mdb_out_7_),
    .Y(_04231_)
  );
  INVX1 _11136_ (
    .A(_00158_),
    .Y(_04232_)
  );
  INVX1 _11137_ (
    .A(eu_mdb_out_8_),
    .Y(_04233_)
  );
  INVX1 _11138_ (
    .A(_00159_),
    .Y(_04234_)
  );
  INVX1 _11139_ (
    .A(eu_mdb_out_9_),
    .Y(_04235_)
  );
  INVX1 _11140_ (
    .A(_00145_),
    .Y(_04236_)
  );
  INVX1 _11141_ (
    .A(eu_mdb_out_10_),
    .Y(_04237_)
  );
  INVX1 _11142_ (
    .A(_00146_),
    .Y(_04238_)
  );
  INVX1 _11143_ (
    .A(eu_mdb_out_11_),
    .Y(_04239_)
  );
  INVX1 _11144_ (
    .A(_00147_),
    .Y(_04240_)
  );
  INVX1 _11145_ (
    .A(eu_mdb_out_12_),
    .Y(_04241_)
  );
  INVX1 _11146_ (
    .A(_00148_),
    .Y(_04242_)
  );
  INVX1 _11147_ (
    .A(eu_mdb_out_13_),
    .Y(_04243_)
  );
  INVX1 _11148_ (
    .A(_00149_),
    .Y(_04244_)
  );
  INVX1 _11149_ (
    .A(eu_mdb_out_14_),
    .Y(_04245_)
  );
  INVX1 _11150_ (
    .A(_00150_),
    .Y(_04246_)
  );
  INVX1 _11151_ (
    .A(eu_mdb_out_15_),
    .Y(_04247_)
  );
  INVX1 _11152_ (
    .A(_00162_),
    .Y(_04165_)
  );
  NAND2X1 _11153_ (
    .A(execution_unit_0.pc_nxt_15_ ),
    .B(fe_mb_en),
    .Y(_04248_)
  );
  INVX1 _11154_ (
    .A(_04248_),
    .Y(mem_backbone_0.fe_pmem_en )
  );
  NAND3X1 _11155_ (
    .A(mem_backbone_0.fe_pmem_en_dly ),
    .B(_04166_),
    .C(_04248_),
    .Y(_04249_)
  );
  MUX2X1 _11156_ (
    .A(mem_backbone_0.pmem_dout_bckup_0_ ),
    .B(pmem_dout_0_),
    .S(_04249_),
    .Y(_04250_)
  );
  INVX1 _11157_ (
    .A(_04250_),
    .Y(_04141_)
  );
  MUX2X1 _11158_ (
    .A(mem_backbone_0.pmem_dout_bckup_1_ ),
    .B(pmem_dout_1_),
    .S(_04249_),
    .Y(_04251_)
  );
  INVX1 _11159_ (
    .A(_04251_),
    .Y(_04148_)
  );
  MUX2X1 _11160_ (
    .A(mem_backbone_0.pmem_dout_bckup_2_ ),
    .B(pmem_dout_2_),
    .S(_04249_),
    .Y(_04252_)
  );
  INVX1 _11161_ (
    .A(_04252_),
    .Y(_04149_)
  );
  MUX2X1 _11162_ (
    .A(mem_backbone_0.pmem_dout_bckup_3_ ),
    .B(pmem_dout_3_),
    .S(_04249_),
    .Y(_04253_)
  );
  INVX1 _11163_ (
    .A(_04253_),
    .Y(_04150_)
  );
  MUX2X1 _11164_ (
    .A(mem_backbone_0.pmem_dout_bckup_4_ ),
    .B(pmem_dout_4_),
    .S(_04249_),
    .Y(_04254_)
  );
  INVX1 _11165_ (
    .A(_04254_),
    .Y(_04151_)
  );
  MUX2X1 _11166_ (
    .A(mem_backbone_0.pmem_dout_bckup_5_ ),
    .B(pmem_dout_5_),
    .S(_04249_),
    .Y(_04255_)
  );
  INVX1 _11167_ (
    .A(_04255_),
    .Y(_04152_)
  );
  MUX2X1 _11168_ (
    .A(mem_backbone_0.pmem_dout_bckup_6_ ),
    .B(pmem_dout_6_),
    .S(_04249_),
    .Y(_04256_)
  );
  INVX1 _11169_ (
    .A(_04256_),
    .Y(_04153_)
  );
  MUX2X1 _11170_ (
    .A(mem_backbone_0.pmem_dout_bckup_7_ ),
    .B(pmem_dout_7_),
    .S(_04249_),
    .Y(_04257_)
  );
  INVX1 _11171_ (
    .A(_04257_),
    .Y(_04154_)
  );
  MUX2X1 _11172_ (
    .A(mem_backbone_0.pmem_dout_bckup_8_ ),
    .B(pmem_dout_8_),
    .S(_04249_),
    .Y(_04258_)
  );
  INVX1 _11173_ (
    .A(_04258_),
    .Y(_04155_)
  );
  MUX2X1 _11174_ (
    .A(_04164_),
    .B(pmem_dout_9_),
    .S(_04249_),
    .Y(_04259_)
  );
  INVX1 _11175_ (
    .A(_04259_),
    .Y(_04156_)
  );
  MUX2X1 _11176_ (
    .A(_04158_),
    .B(pmem_dout_10_),
    .S(_04249_),
    .Y(_04260_)
  );
  INVX1 _11177_ (
    .A(_04260_),
    .Y(_04142_)
  );
  MUX2X1 _11178_ (
    .A(_04159_),
    .B(pmem_dout_11_),
    .S(_04249_),
    .Y(_04261_)
  );
  INVX1 _11179_ (
    .A(_04261_),
    .Y(_04143_)
  );
  MUX2X1 _11180_ (
    .A(_04160_),
    .B(pmem_dout_12_),
    .S(_04249_),
    .Y(_04262_)
  );
  INVX1 _11181_ (
    .A(_04262_),
    .Y(_04144_)
  );
  MUX2X1 _11182_ (
    .A(_04161_),
    .B(pmem_dout_13_),
    .S(_04249_),
    .Y(_04263_)
  );
  INVX1 _11183_ (
    .A(_04263_),
    .Y(_04145_)
  );
  MUX2X1 _11184_ (
    .A(_04162_),
    .B(pmem_dout_14_),
    .S(_04249_),
    .Y(_04264_)
  );
  INVX1 _11185_ (
    .A(_04264_),
    .Y(_04146_)
  );
  MUX2X1 _11186_ (
    .A(_04163_),
    .B(pmem_dout_15_),
    .S(_04249_),
    .Y(_04265_)
  );
  INVX1 _11187_ (
    .A(_04265_),
    .Y(_04147_)
  );
  NOR2X1 _11188_ (
    .A(_04200_),
    .B(dbg_0.UNUSED_eu_mab_15_ ),
    .Y(_04266_)
  );
  INVX1 _11189_ (
    .A(_04266_),
    .Y(_04267_)
  );
  NAND3X1 _11190_ (
    .A(_04185_),
    .B(dbg_0.dbg_mem_addr_14_ ),
    .C(dbg_0.dbg_mem_en ),
    .Y(_04268_)
  );
  INVX1 _11191_ (
    .A(_04268_),
    .Y(_04269_)
  );
  AOI21X1 _11192_ (
    .A(dbg_0.UNUSED_eu_mab_14_ ),
    .B(_04266_),
    .C(_04268_),
    .Y(_04270_)
  );
  MUX2X1 _11193_ (
    .A(dbg_0.dbg_mem_wr_0_ ),
    .B(dbg_0.UNUSED_eu_mb_wr_0_ ),
    .S(_04270_),
    .Y(_00081_)
  );
  MUX2X1 _11194_ (
    .A(dbg_0.dbg_mem_wr_1_ ),
    .B(dbg_0.UNUSED_eu_mb_wr_1_ ),
    .S(_04270_),
    .Y(_00082_)
  );
  MUX2X1 _11195_ (
    .A(_04199_),
    .B(_04213_),
    .S(_04270_),
    .Y(_00051_)
  );
  MUX2X1 _11196_ (
    .A(_04198_),
    .B(_04212_),
    .S(_04270_),
    .Y(_00055_)
  );
  MUX2X1 _11197_ (
    .A(_04197_),
    .B(_04211_),
    .S(_04270_),
    .Y(_00056_)
  );
  MUX2X1 _11198_ (
    .A(_04196_),
    .B(_04210_),
    .S(_04270_),
    .Y(_00057_)
  );
  MUX2X1 _11199_ (
    .A(_04195_),
    .B(_04209_),
    .S(_04270_),
    .Y(_00058_)
  );
  MUX2X1 _11200_ (
    .A(_04194_),
    .B(_04208_),
    .S(_04270_),
    .Y(_00059_)
  );
  MUX2X1 _11201_ (
    .A(_04193_),
    .B(_04207_),
    .S(_04270_),
    .Y(_00060_)
  );
  MUX2X1 _11202_ (
    .A(_04192_),
    .B(_04206_),
    .S(_04270_),
    .Y(_00061_)
  );
  MUX2X1 _11203_ (
    .A(_04191_),
    .B(_04205_),
    .S(_04270_),
    .Y(_00062_)
  );
  MUX2X1 _11204_ (
    .A(_04190_),
    .B(_04204_),
    .S(_04270_),
    .Y(_00063_)
  );
  MUX2X1 _11205_ (
    .A(_04189_),
    .B(_04203_),
    .S(_04270_),
    .Y(_00052_)
  );
  MUX2X1 _11206_ (
    .A(_04188_),
    .B(_04202_),
    .S(_04270_),
    .Y(_00053_)
  );
  MUX2X1 _11207_ (
    .A(_04187_),
    .B(_04201_),
    .S(_04270_),
    .Y(_00054_)
  );
  MUX2X1 _11208_ (
    .A(_04216_),
    .B(_04217_),
    .S(_04270_),
    .Y(_00065_)
  );
  MUX2X1 _11209_ (
    .A(_04218_),
    .B(_04219_),
    .S(_04270_),
    .Y(_00072_)
  );
  MUX2X1 _11210_ (
    .A(_04220_),
    .B(_04221_),
    .S(_04270_),
    .Y(_00073_)
  );
  MUX2X1 _11211_ (
    .A(_04222_),
    .B(_04223_),
    .S(_04270_),
    .Y(_00074_)
  );
  MUX2X1 _11212_ (
    .A(_04224_),
    .B(_04225_),
    .S(_04270_),
    .Y(_00075_)
  );
  MUX2X1 _11213_ (
    .A(_04226_),
    .B(_04227_),
    .S(_04270_),
    .Y(_00076_)
  );
  MUX2X1 _11214_ (
    .A(_04228_),
    .B(_04229_),
    .S(_04270_),
    .Y(_00077_)
  );
  MUX2X1 _11215_ (
    .A(_04230_),
    .B(_04231_),
    .S(_04270_),
    .Y(_00078_)
  );
  MUX2X1 _11216_ (
    .A(_04232_),
    .B(_04233_),
    .S(_04270_),
    .Y(_00079_)
  );
  MUX2X1 _11217_ (
    .A(_04234_),
    .B(_04235_),
    .S(_04270_),
    .Y(_00080_)
  );
  MUX2X1 _11218_ (
    .A(_04236_),
    .B(_04237_),
    .S(_04270_),
    .Y(_00066_)
  );
  MUX2X1 _11219_ (
    .A(_04238_),
    .B(_04239_),
    .S(_04270_),
    .Y(_00067_)
  );
  MUX2X1 _11220_ (
    .A(_04240_),
    .B(_04241_),
    .S(_04270_),
    .Y(_00068_)
  );
  MUX2X1 _11221_ (
    .A(_04242_),
    .B(_04243_),
    .S(_04270_),
    .Y(_00069_)
  );
  MUX2X1 _11222_ (
    .A(_04244_),
    .B(_04245_),
    .S(_04270_),
    .Y(_00070_)
  );
  MUX2X1 _11223_ (
    .A(_04246_),
    .B(_04247_),
    .S(_04270_),
    .Y(_00071_)
  );
  OR2X1 _11224_ (
    .A(dbg_0.UNUSED_eu_mb_wr_0_ ),
    .B(dbg_0.UNUSED_eu_mb_wr_1_ ),
    .Y(_04271_)
  );
  NAND2X1 _11225_ (
    .A(dbg_0.UNUSED_eu_mb_en ),
    .B(dbg_0.UNUSED_eu_mab_15_ ),
    .Y(_04272_)
  );
  OR2X1 _11226_ (
    .A(_04271_),
    .B(_04272_),
    .Y(_04273_)
  );
  INVX1 _11227_ (
    .A(_04273_),
    .Y(mem_backbone_0.eu_pmem_en )
  );
  OAI21X1 _11228_ (
    .A(_04271_),
    .B(_04272_),
    .C(_04248_),
    .Y(_04274_)
  );
  NAND2X1 _11229_ (
    .A(dbg_0.dbg_mem_addr_15_ ),
    .B(dbg_0.dbg_mem_en ),
    .Y(_04275_)
  );
  NOR2X1 _11230_ (
    .A(_04274_),
    .B(_04275_),
    .Y(mem_backbone_0.ext_pmem_en )
  );
  NAND2X1 _11231_ (
    .A(dbg_0.dbg_mem_wr_0_ ),
    .B(mem_backbone_0.ext_pmem_en ),
    .Y(_00160_)
  );
  NAND2X1 _11232_ (
    .A(dbg_0.dbg_mem_wr_1_ ),
    .B(mem_backbone_0.ext_pmem_en ),
    .Y(_00161_)
  );
  MUX2X1 _11233_ (
    .A(execution_unit_0.pc_nxt_1_ ),
    .B(dbg_0.UNUSED_eu_mab_1_ ),
    .S(_04273_),
    .Y(_04276_)
  );
  MUX2X1 _11234_ (
    .A(_04199_),
    .B(_04276_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00129_)
  );
  MUX2X1 _11235_ (
    .A(execution_unit_0.pc_nxt_2_ ),
    .B(dbg_0.UNUSED_eu_mab_2_ ),
    .S(_04273_),
    .Y(_04277_)
  );
  MUX2X1 _11236_ (
    .A(_04198_),
    .B(_04277_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00134_)
  );
  MUX2X1 _11237_ (
    .A(execution_unit_0.pc_nxt_3_ ),
    .B(dbg_0.UNUSED_eu_mab_3_ ),
    .S(_04273_),
    .Y(_04278_)
  );
  MUX2X1 _11238_ (
    .A(_04197_),
    .B(_04278_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00135_)
  );
  MUX2X1 _11239_ (
    .A(execution_unit_0.pc_nxt_4_ ),
    .B(dbg_0.UNUSED_eu_mab_4_ ),
    .S(_04273_),
    .Y(_04279_)
  );
  MUX2X1 _11240_ (
    .A(_04196_),
    .B(_04279_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00136_)
  );
  MUX2X1 _11241_ (
    .A(execution_unit_0.pc_nxt_5_ ),
    .B(dbg_0.UNUSED_eu_mab_5_ ),
    .S(_04273_),
    .Y(_04280_)
  );
  MUX2X1 _11242_ (
    .A(_04195_),
    .B(_04280_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00137_)
  );
  MUX2X1 _11243_ (
    .A(execution_unit_0.pc_nxt_6_ ),
    .B(dbg_0.UNUSED_eu_mab_6_ ),
    .S(_04273_),
    .Y(_04281_)
  );
  MUX2X1 _11244_ (
    .A(_04194_),
    .B(_04281_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00138_)
  );
  MUX2X1 _11245_ (
    .A(execution_unit_0.pc_nxt_7_ ),
    .B(dbg_0.UNUSED_eu_mab_7_ ),
    .S(_04273_),
    .Y(_04282_)
  );
  MUX2X1 _11246_ (
    .A(_04193_),
    .B(_04282_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00139_)
  );
  MUX2X1 _11247_ (
    .A(execution_unit_0.pc_nxt_8_ ),
    .B(dbg_0.UNUSED_eu_mab_8_ ),
    .S(_04273_),
    .Y(_04283_)
  );
  MUX2X1 _11248_ (
    .A(_04192_),
    .B(_04283_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00140_)
  );
  MUX2X1 _11249_ (
    .A(execution_unit_0.pc_nxt_9_ ),
    .B(dbg_0.UNUSED_eu_mab_9_ ),
    .S(_04273_),
    .Y(_04284_)
  );
  MUX2X1 _11250_ (
    .A(_04191_),
    .B(_04284_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00141_)
  );
  MUX2X1 _11251_ (
    .A(execution_unit_0.pc_nxt_10_ ),
    .B(dbg_0.UNUSED_eu_mab_10_ ),
    .S(_04273_),
    .Y(_04285_)
  );
  MUX2X1 _11252_ (
    .A(_04190_),
    .B(_04285_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00142_)
  );
  MUX2X1 _11253_ (
    .A(execution_unit_0.pc_nxt_11_ ),
    .B(dbg_0.UNUSED_eu_mab_11_ ),
    .S(_04273_),
    .Y(_04286_)
  );
  MUX2X1 _11254_ (
    .A(_04189_),
    .B(_04286_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00130_)
  );
  MUX2X1 _11255_ (
    .A(execution_unit_0.pc_nxt_12_ ),
    .B(dbg_0.UNUSED_eu_mab_12_ ),
    .S(_04273_),
    .Y(_04287_)
  );
  MUX2X1 _11256_ (
    .A(_04188_),
    .B(_04287_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00131_)
  );
  MUX2X1 _11257_ (
    .A(execution_unit_0.pc_nxt_13_ ),
    .B(dbg_0.UNUSED_eu_mab_13_ ),
    .S(_04273_),
    .Y(_04288_)
  );
  MUX2X1 _11258_ (
    .A(_04187_),
    .B(_04288_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00132_)
  );
  MUX2X1 _11259_ (
    .A(execution_unit_0.pc_nxt_14_ ),
    .B(dbg_0.UNUSED_eu_mab_14_ ),
    .S(_04273_),
    .Y(_04289_)
  );
  MUX2X1 _11260_ (
    .A(_04186_),
    .B(_04289_),
    .S(mem_backbone_0.ext_pmem_en ),
    .Y(_00133_)
  );
  NOR3X1 _11261_ (
    .A(_04200_),
    .B(dbg_0.UNUSED_eu_mab_15_ ),
    .C(dbg_0.UNUSED_eu_mab_14_ ),
    .Y(mem_backbone_0.eu_per_en )
  );
  NAND3X1 _11262_ (
    .A(_04185_),
    .B(_04186_),
    .C(dbg_0.dbg_mem_en ),
    .Y(_04290_)
  );
  NOR2X1 _11263_ (
    .A(mem_backbone_0.eu_per_en ),
    .B(_04290_),
    .Y(mem_backbone_0.ext_per_en )
  );
  MUX2X1 _11264_ (
    .A(_04184_),
    .B(_04183_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00127_)
  );
  MUX2X1 _11265_ (
    .A(_04215_),
    .B(_04214_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00128_)
  );
  MUX2X1 _11266_ (
    .A(_04199_),
    .B(_04213_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00097_)
  );
  MUX2X1 _11267_ (
    .A(_04198_),
    .B(_04212_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00101_)
  );
  MUX2X1 _11268_ (
    .A(_04197_),
    .B(_04211_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00102_)
  );
  MUX2X1 _11269_ (
    .A(_04196_),
    .B(_04210_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00103_)
  );
  MUX2X1 _11270_ (
    .A(_04195_),
    .B(_04209_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00104_)
  );
  MUX2X1 _11271_ (
    .A(_04194_),
    .B(_04208_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00105_)
  );
  MUX2X1 _11272_ (
    .A(_04193_),
    .B(_04207_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00106_)
  );
  MUX2X1 _11273_ (
    .A(_04192_),
    .B(_04206_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00107_)
  );
  MUX2X1 _11274_ (
    .A(_04191_),
    .B(_04205_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00108_)
  );
  MUX2X1 _11275_ (
    .A(_04190_),
    .B(_04204_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00109_)
  );
  MUX2X1 _11276_ (
    .A(_04189_),
    .B(_04203_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00098_)
  );
  MUX2X1 _11277_ (
    .A(_04188_),
    .B(_04202_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00099_)
  );
  MUX2X1 _11278_ (
    .A(_04187_),
    .B(_04201_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00100_)
  );
  MUX2X1 _11279_ (
    .A(_04216_),
    .B(_04217_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00110_)
  );
  MUX2X1 _11280_ (
    .A(_04218_),
    .B(_04219_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00117_)
  );
  MUX2X1 _11281_ (
    .A(_04220_),
    .B(_04221_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00118_)
  );
  MUX2X1 _11282_ (
    .A(_04222_),
    .B(_04223_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00119_)
  );
  MUX2X1 _11283_ (
    .A(_04224_),
    .B(_04225_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00120_)
  );
  MUX2X1 _11284_ (
    .A(_04226_),
    .B(_04227_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00121_)
  );
  MUX2X1 _11285_ (
    .A(_04228_),
    .B(_04229_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00122_)
  );
  MUX2X1 _11286_ (
    .A(_04230_),
    .B(_04231_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00123_)
  );
  MUX2X1 _11287_ (
    .A(_04232_),
    .B(_04233_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00124_)
  );
  MUX2X1 _11288_ (
    .A(_04234_),
    .B(_04235_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00125_)
  );
  MUX2X1 _11289_ (
    .A(_04236_),
    .B(_04237_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00111_)
  );
  MUX2X1 _11290_ (
    .A(_04238_),
    .B(_04239_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00112_)
  );
  MUX2X1 _11291_ (
    .A(_04240_),
    .B(_04241_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00113_)
  );
  MUX2X1 _11292_ (
    .A(_04242_),
    .B(_04243_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00114_)
  );
  MUX2X1 _11293_ (
    .A(_04244_),
    .B(_04245_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00115_)
  );
  MUX2X1 _11294_ (
    .A(_04246_),
    .B(_04247_),
    .S(mem_backbone_0.ext_per_en ),
    .Y(_00116_)
  );
  NAND2X1 _11295_ (
    .A(mem_backbone_0.pmem_dout_bckup_0_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04291_)
  );
  OAI21X1 _11296_ (
    .A(_04167_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04291_),
    .Y(dbg_0.fe_mdb_in_0_ )
  );
  NAND2X1 _11297_ (
    .A(mem_backbone_0.pmem_dout_bckup_1_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04292_)
  );
  OAI21X1 _11298_ (
    .A(_04168_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04292_),
    .Y(dbg_0.fe_mdb_in_1_ )
  );
  NAND2X1 _11299_ (
    .A(mem_backbone_0.pmem_dout_bckup_2_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04293_)
  );
  OAI21X1 _11300_ (
    .A(_04169_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04293_),
    .Y(dbg_0.fe_mdb_in_2_ )
  );
  NAND2X1 _11301_ (
    .A(mem_backbone_0.pmem_dout_bckup_3_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04294_)
  );
  OAI21X1 _11302_ (
    .A(_04170_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04294_),
    .Y(dbg_0.fe_mdb_in_3_ )
  );
  NAND2X1 _11303_ (
    .A(mem_backbone_0.pmem_dout_bckup_4_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04295_)
  );
  OAI21X1 _11304_ (
    .A(_04171_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04295_),
    .Y(dbg_0.fe_mdb_in_4_ )
  );
  NAND2X1 _11305_ (
    .A(mem_backbone_0.pmem_dout_bckup_5_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04296_)
  );
  OAI21X1 _11306_ (
    .A(_04172_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04296_),
    .Y(dbg_0.fe_mdb_in_5_ )
  );
  NAND2X1 _11307_ (
    .A(mem_backbone_0.pmem_dout_bckup_6_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04297_)
  );
  OAI21X1 _11308_ (
    .A(_04173_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04297_),
    .Y(dbg_0.fe_mdb_in_6_ )
  );
  NAND2X1 _11309_ (
    .A(mem_backbone_0.pmem_dout_bckup_7_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04298_)
  );
  OAI21X1 _11310_ (
    .A(_04174_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04298_),
    .Y(dbg_0.fe_mdb_in_7_ )
  );
  NAND2X1 _11311_ (
    .A(mem_backbone_0.pmem_dout_bckup_8_ ),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04299_)
  );
  OAI21X1 _11312_ (
    .A(_04175_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04299_),
    .Y(dbg_0.fe_mdb_in_8_ )
  );
  NAND2X1 _11313_ (
    .A(_04164_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04300_)
  );
  OAI21X1 _11314_ (
    .A(_04176_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04300_),
    .Y(dbg_0.fe_mdb_in_9_ )
  );
  NAND2X1 _11315_ (
    .A(_04158_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04301_)
  );
  OAI21X1 _11316_ (
    .A(_04177_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04301_),
    .Y(dbg_0.fe_mdb_in_10_ )
  );
  NAND2X1 _11317_ (
    .A(_04159_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04302_)
  );
  OAI21X1 _11318_ (
    .A(_04178_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04302_),
    .Y(dbg_0.fe_mdb_in_11_ )
  );
  NAND2X1 _11319_ (
    .A(_04160_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04303_)
  );
  OAI21X1 _11320_ (
    .A(_04179_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04303_),
    .Y(dbg_0.fe_mdb_in_12_ )
  );
  NAND2X1 _11321_ (
    .A(_04161_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04304_)
  );
  OAI21X1 _11322_ (
    .A(_04180_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04304_),
    .Y(dbg_0.fe_mdb_in_13_ )
  );
  NAND2X1 _11323_ (
    .A(_04162_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04305_)
  );
  OAI21X1 _11324_ (
    .A(_04181_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04305_),
    .Y(dbg_0.fe_mdb_in_14_ )
  );
  NAND2X1 _11325_ (
    .A(_04163_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04306_)
  );
  OAI21X1 _11326_ (
    .A(_04182_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .C(_04306_),
    .Y(dbg_0.fe_mdb_in_15_ )
  );
  MUX2X1 _11327_ (
    .A(mem_backbone_0.per_dout_val_0_ ),
    .B(dmem_dout_0_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04307_)
  );
  NAND2X1 _11328_ (
    .A(pmem_dout_0_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04308_)
  );
  OAI21X1 _11329_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04307_),
    .C(_04308_),
    .Y(eu_mdb_in_0_)
  );
  MUX2X1 _11330_ (
    .A(mem_backbone_0.per_dout_val_1_ ),
    .B(dmem_dout_1_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04309_)
  );
  NAND2X1 _11331_ (
    .A(pmem_dout_1_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04310_)
  );
  OAI21X1 _11332_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04309_),
    .C(_04310_),
    .Y(eu_mdb_in_1_)
  );
  MUX2X1 _11333_ (
    .A(mem_backbone_0.per_dout_val_2_ ),
    .B(dmem_dout_2_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04311_)
  );
  NAND2X1 _11334_ (
    .A(pmem_dout_2_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04312_)
  );
  OAI21X1 _11335_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04311_),
    .C(_04312_),
    .Y(eu_mdb_in_2_)
  );
  MUX2X1 _11336_ (
    .A(mem_backbone_0.per_dout_val_3_ ),
    .B(dmem_dout_3_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04313_)
  );
  NAND2X1 _11337_ (
    .A(pmem_dout_3_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04314_)
  );
  OAI21X1 _11338_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04313_),
    .C(_04314_),
    .Y(eu_mdb_in_3_)
  );
  MUX2X1 _11339_ (
    .A(mem_backbone_0.per_dout_val_4_ ),
    .B(dmem_dout_4_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04315_)
  );
  NAND2X1 _11340_ (
    .A(pmem_dout_4_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04316_)
  );
  OAI21X1 _11341_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04315_),
    .C(_04316_),
    .Y(eu_mdb_in_4_)
  );
  MUX2X1 _11342_ (
    .A(mem_backbone_0.per_dout_val_5_ ),
    .B(dmem_dout_5_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04317_)
  );
  NAND2X1 _11343_ (
    .A(pmem_dout_5_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04318_)
  );
  OAI21X1 _11344_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04317_),
    .C(_04318_),
    .Y(eu_mdb_in_5_)
  );
  MUX2X1 _11345_ (
    .A(mem_backbone_0.per_dout_val_6_ ),
    .B(dmem_dout_6_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04319_)
  );
  NAND2X1 _11346_ (
    .A(pmem_dout_6_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04320_)
  );
  OAI21X1 _11347_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04319_),
    .C(_04320_),
    .Y(eu_mdb_in_6_)
  );
  MUX2X1 _11348_ (
    .A(mem_backbone_0.per_dout_val_7_ ),
    .B(dmem_dout_7_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04321_)
  );
  NAND2X1 _11349_ (
    .A(pmem_dout_7_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04322_)
  );
  OAI21X1 _11350_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04321_),
    .C(_04322_),
    .Y(eu_mdb_in_7_)
  );
  MUX2X1 _11351_ (
    .A(mem_backbone_0.per_dout_val_8_ ),
    .B(dmem_dout_8_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04323_)
  );
  NAND2X1 _11352_ (
    .A(pmem_dout_8_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04324_)
  );
  OAI21X1 _11353_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04323_),
    .C(_04324_),
    .Y(eu_mdb_in_8_)
  );
  MUX2X1 _11354_ (
    .A(mem_backbone_0.per_dout_val_9_ ),
    .B(dmem_dout_9_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04325_)
  );
  NAND2X1 _11355_ (
    .A(pmem_dout_9_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04326_)
  );
  OAI21X1 _11356_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04325_),
    .C(_04326_),
    .Y(eu_mdb_in_9_)
  );
  MUX2X1 _11357_ (
    .A(mem_backbone_0.per_dout_val_10_ ),
    .B(dmem_dout_10_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04327_)
  );
  NAND2X1 _11358_ (
    .A(pmem_dout_10_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04328_)
  );
  OAI21X1 _11359_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04327_),
    .C(_04328_),
    .Y(eu_mdb_in_10_)
  );
  MUX2X1 _11360_ (
    .A(mem_backbone_0.per_dout_val_11_ ),
    .B(dmem_dout_11_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04329_)
  );
  NAND2X1 _11361_ (
    .A(pmem_dout_11_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04330_)
  );
  OAI21X1 _11362_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04329_),
    .C(_04330_),
    .Y(eu_mdb_in_11_)
  );
  MUX2X1 _11363_ (
    .A(mem_backbone_0.per_dout_val_12_ ),
    .B(dmem_dout_12_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04331_)
  );
  NAND2X1 _11364_ (
    .A(pmem_dout_12_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04332_)
  );
  OAI21X1 _11365_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04331_),
    .C(_04332_),
    .Y(eu_mdb_in_12_)
  );
  MUX2X1 _11366_ (
    .A(mem_backbone_0.per_dout_val_13_ ),
    .B(dmem_dout_13_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04333_)
  );
  NAND2X1 _11367_ (
    .A(pmem_dout_13_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04334_)
  );
  OAI21X1 _11368_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04333_),
    .C(_04334_),
    .Y(eu_mdb_in_13_)
  );
  MUX2X1 _11369_ (
    .A(mem_backbone_0.per_dout_val_14_ ),
    .B(dmem_dout_14_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04335_)
  );
  NAND2X1 _11370_ (
    .A(pmem_dout_14_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04336_)
  );
  OAI21X1 _11371_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04335_),
    .C(_04336_),
    .Y(eu_mdb_in_14_)
  );
  MUX2X1 _11372_ (
    .A(mem_backbone_0.per_dout_val_15_ ),
    .B(dmem_dout_15_),
    .S(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .Y(_04337_)
  );
  NAND2X1 _11373_ (
    .A(pmem_dout_15_),
    .B(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .Y(_04338_)
  );
  OAI21X1 _11374_ (
    .A(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .B(_04337_),
    .C(_04338_),
    .Y(eu_mdb_in_15_)
  );
  MUX2X1 _11375_ (
    .A(mem_backbone_0.per_dout_val_0_ ),
    .B(dmem_dout_0_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04339_)
  );
  NAND2X1 _11376_ (
    .A(pmem_dout_0_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04340_)
  );
  OAI21X1 _11377_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04339_),
    .C(_04340_),
    .Y(dbg_0.dbg_mem_din_0_ )
  );
  MUX2X1 _11378_ (
    .A(mem_backbone_0.per_dout_val_1_ ),
    .B(dmem_dout_1_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04341_)
  );
  NAND2X1 _11379_ (
    .A(pmem_dout_1_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04342_)
  );
  OAI21X1 _11380_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04341_),
    .C(_04342_),
    .Y(dbg_0.dbg_mem_din_1_ )
  );
  MUX2X1 _11381_ (
    .A(mem_backbone_0.per_dout_val_2_ ),
    .B(dmem_dout_2_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04343_)
  );
  NAND2X1 _11382_ (
    .A(pmem_dout_2_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04344_)
  );
  OAI21X1 _11383_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04343_),
    .C(_04344_),
    .Y(dbg_0.dbg_mem_din_2_ )
  );
  MUX2X1 _11384_ (
    .A(mem_backbone_0.per_dout_val_3_ ),
    .B(dmem_dout_3_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04345_)
  );
  NAND2X1 _11385_ (
    .A(pmem_dout_3_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04346_)
  );
  OAI21X1 _11386_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04345_),
    .C(_04346_),
    .Y(dbg_0.dbg_mem_din_3_ )
  );
  MUX2X1 _11387_ (
    .A(mem_backbone_0.per_dout_val_4_ ),
    .B(dmem_dout_4_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04347_)
  );
  NAND2X1 _11388_ (
    .A(pmem_dout_4_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04348_)
  );
  OAI21X1 _11389_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04347_),
    .C(_04348_),
    .Y(dbg_0.dbg_mem_din_4_ )
  );
  MUX2X1 _11390_ (
    .A(mem_backbone_0.per_dout_val_5_ ),
    .B(dmem_dout_5_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04349_)
  );
  NAND2X1 _11391_ (
    .A(pmem_dout_5_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04350_)
  );
  OAI21X1 _11392_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04349_),
    .C(_04350_),
    .Y(dbg_0.dbg_mem_din_5_ )
  );
  MUX2X1 _11393_ (
    .A(mem_backbone_0.per_dout_val_6_ ),
    .B(dmem_dout_6_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04351_)
  );
  NAND2X1 _11394_ (
    .A(pmem_dout_6_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04352_)
  );
  OAI21X1 _11395_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04351_),
    .C(_04352_),
    .Y(dbg_0.dbg_mem_din_6_ )
  );
  MUX2X1 _11396_ (
    .A(mem_backbone_0.per_dout_val_7_ ),
    .B(dmem_dout_7_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04353_)
  );
  NAND2X1 _11397_ (
    .A(pmem_dout_7_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04354_)
  );
  OAI21X1 _11398_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04353_),
    .C(_04354_),
    .Y(dbg_0.dbg_mem_din_7_ )
  );
  MUX2X1 _11399_ (
    .A(mem_backbone_0.per_dout_val_8_ ),
    .B(dmem_dout_8_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04355_)
  );
  NAND2X1 _11400_ (
    .A(pmem_dout_8_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04356_)
  );
  OAI21X1 _11401_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04355_),
    .C(_04356_),
    .Y(dbg_0.dbg_mem_din_8_ )
  );
  MUX2X1 _11402_ (
    .A(mem_backbone_0.per_dout_val_9_ ),
    .B(dmem_dout_9_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04357_)
  );
  NAND2X1 _11403_ (
    .A(pmem_dout_9_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04358_)
  );
  OAI21X1 _11404_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04357_),
    .C(_04358_),
    .Y(dbg_0.dbg_mem_din_9_ )
  );
  MUX2X1 _11405_ (
    .A(mem_backbone_0.per_dout_val_10_ ),
    .B(dmem_dout_10_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04359_)
  );
  NAND2X1 _11406_ (
    .A(pmem_dout_10_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04360_)
  );
  OAI21X1 _11407_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04359_),
    .C(_04360_),
    .Y(dbg_0.dbg_mem_din_10_ )
  );
  MUX2X1 _11408_ (
    .A(mem_backbone_0.per_dout_val_11_ ),
    .B(dmem_dout_11_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04361_)
  );
  NAND2X1 _11409_ (
    .A(pmem_dout_11_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04362_)
  );
  OAI21X1 _11410_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04361_),
    .C(_04362_),
    .Y(dbg_0.dbg_mem_din_11_ )
  );
  MUX2X1 _11411_ (
    .A(mem_backbone_0.per_dout_val_12_ ),
    .B(dmem_dout_12_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04363_)
  );
  NAND2X1 _11412_ (
    .A(pmem_dout_12_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04364_)
  );
  OAI21X1 _11413_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04363_),
    .C(_04364_),
    .Y(dbg_0.dbg_mem_din_12_ )
  );
  MUX2X1 _11414_ (
    .A(mem_backbone_0.per_dout_val_13_ ),
    .B(dmem_dout_13_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04365_)
  );
  NAND2X1 _11415_ (
    .A(pmem_dout_13_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04366_)
  );
  OAI21X1 _11416_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04365_),
    .C(_04366_),
    .Y(dbg_0.dbg_mem_din_13_ )
  );
  MUX2X1 _11417_ (
    .A(mem_backbone_0.per_dout_val_14_ ),
    .B(dmem_dout_14_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04367_)
  );
  NAND2X1 _11418_ (
    .A(pmem_dout_14_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04368_)
  );
  OAI21X1 _11419_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04367_),
    .C(_04368_),
    .Y(dbg_0.dbg_mem_din_14_ )
  );
  MUX2X1 _11420_ (
    .A(mem_backbone_0.per_dout_val_15_ ),
    .B(dmem_dout_15_),
    .S(mem_backbone_0.ext_mem_din_sel_0_ ),
    .Y(_04369_)
  );
  NAND2X1 _11421_ (
    .A(pmem_dout_15_),
    .B(mem_backbone_0.ext_mem_din_sel_1_ ),
    .Y(_04370_)
  );
  OAI21X1 _11422_ (
    .A(mem_backbone_0.ext_mem_din_sel_1_ ),
    .B(_04369_),
    .C(_04370_),
    .Y(dbg_0.dbg_mem_din_15_ )
  );
  AOI21X1 _11423_ (
    .A(dbg_0.UNUSED_eu_mab_14_ ),
    .B(_04266_),
    .C(_04269_),
    .Y(_00064_)
  );
  NOR2X1 _11424_ (
    .A(_04274_),
    .B(mem_backbone_0.ext_pmem_en ),
    .Y(_00143_)
  );
  NOR2X1 _11425_ (
    .A(mem_backbone_0.fe_pmem_en_dly ),
    .B(_04248_),
    .Y(_04371_)
  );
  NAND2X1 _11426_ (
    .A(_04166_),
    .B(mem_backbone_0.pmem_dout_bckup_sel ),
    .Y(_04372_)
  );
  OAI21X1 _11427_ (
    .A(_04371_),
    .B(_04372_),
    .C(_04249_),
    .Y(_04157_)
  );
  NOR2X1 _11428_ (
    .A(_04248_),
    .B(_04273_),
    .Y(fe_pmem_wait)
  );
  OAI21X1 _11429_ (
    .A(dbg_0.UNUSED_eu_mab_14_ ),
    .B(_04267_),
    .C(_04290_),
    .Y(_00126_)
  );
  DFFSR _11430_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.ext_per_en ),
    .Q(mem_backbone_0.ext_mem_din_sel_0_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11431_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.ext_pmem_en ),
    .Q(mem_backbone_0.ext_mem_din_sel_1_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11432_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.eu_per_en ),
    .Q(mem_backbone_0.eu_mdb_in_sel_0_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11433_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.eu_pmem_en ),
    .Q(mem_backbone_0.eu_mdb_in_sel_1_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11434_ (
    .CLK(dco_clk),
    .D(_04157_),
    .Q(mem_backbone_0.pmem_dout_bckup_sel ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11435_ (
    .CLK(dco_clk),
    .D(_04141_),
    .Q(mem_backbone_0.pmem_dout_bckup_0_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11436_ (
    .CLK(dco_clk),
    .D(_04148_),
    .Q(mem_backbone_0.pmem_dout_bckup_1_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11437_ (
    .CLK(dco_clk),
    .D(_04149_),
    .Q(mem_backbone_0.pmem_dout_bckup_2_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11438_ (
    .CLK(dco_clk),
    .D(_04150_),
    .Q(mem_backbone_0.pmem_dout_bckup_3_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11439_ (
    .CLK(dco_clk),
    .D(_04151_),
    .Q(mem_backbone_0.pmem_dout_bckup_4_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11440_ (
    .CLK(dco_clk),
    .D(_04152_),
    .Q(mem_backbone_0.pmem_dout_bckup_5_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11441_ (
    .CLK(dco_clk),
    .D(_04153_),
    .Q(mem_backbone_0.pmem_dout_bckup_6_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11442_ (
    .CLK(dco_clk),
    .D(_04154_),
    .Q(mem_backbone_0.pmem_dout_bckup_7_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11443_ (
    .CLK(dco_clk),
    .D(_04155_),
    .Q(mem_backbone_0.pmem_dout_bckup_8_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11444_ (
    .CLK(dco_clk),
    .D(_04156_),
    .Q(_04164_),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11445_ (
    .CLK(dco_clk),
    .D(_04142_),
    .Q(_04158_),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11446_ (
    .CLK(dco_clk),
    .D(_04143_),
    .Q(_04159_),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11447_ (
    .CLK(dco_clk),
    .D(_04144_),
    .Q(_04160_),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11448_ (
    .CLK(dco_clk),
    .D(_04145_),
    .Q(_04161_),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11449_ (
    .CLK(dco_clk),
    .D(_04146_),
    .Q(_04162_),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11450_ (
    .CLK(dco_clk),
    .D(_04147_),
    .Q(_04163_),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11451_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.fe_pmem_en ),
    .Q(mem_backbone_0.fe_pmem_en_dly ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11452_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_0_ ),
    .Q(mem_backbone_0.per_dout_val_0_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11453_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_1_ ),
    .Q(mem_backbone_0.per_dout_val_1_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11454_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_2_ ),
    .Q(mem_backbone_0.per_dout_val_2_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11455_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_3_ ),
    .Q(mem_backbone_0.per_dout_val_3_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11456_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_4_ ),
    .Q(mem_backbone_0.per_dout_val_4_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11457_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_5_ ),
    .Q(mem_backbone_0.per_dout_val_5_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11458_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_6_ ),
    .Q(mem_backbone_0.per_dout_val_6_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11459_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_7_ ),
    .Q(mem_backbone_0.per_dout_val_7_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11460_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_8_ ),
    .Q(mem_backbone_0.per_dout_val_8_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11461_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_9_ ),
    .Q(mem_backbone_0.per_dout_val_9_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11462_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_10_ ),
    .Q(mem_backbone_0.per_dout_val_10_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11463_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_11_ ),
    .Q(mem_backbone_0.per_dout_val_11_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11464_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_12_ ),
    .Q(mem_backbone_0.per_dout_val_12_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11465_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_13_ ),
    .Q(mem_backbone_0.per_dout_val_13_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11466_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_14_ ),
    .Q(mem_backbone_0.per_dout_val_14_ ),
    .R(_04165_),
    .S(1'h1)
  );
  DFFSR _11467_ (
    .CLK(dco_clk),
    .D(mem_backbone_0.per_dout_15_ ),
    .Q(mem_backbone_0.per_dout_val_15_ ),
    .R(_04165_),
    .S(1'h1)
  );
  INVX1 _11468_ (
    .A(_00097_),
    .Y(_05042_)
  );
  INVX1 _11469_ (
    .A(_00104_),
    .Y(_05043_)
  );
  INVX1 _11470_ (
    .A(_00106_),
    .Y(_05044_)
  );
  INVX1 _11471_ (
    .A(_00107_),
    .Y(_05045_)
  );
  INVX1 _11472_ (
    .A(_00100_),
    .Y(_05046_)
  );
  INVX1 _11473_ (
    .A(multiplier_0.cycle_0_ ),
    .Y(_05047_)
  );
  INVX1 _11474_ (
    .A(multiplier_0.cycle_1_ ),
    .Y(_05048_)
  );
  INVX1 _11475_ (
    .A(multiplier_0.sign_sel ),
    .Y(_05049_)
  );
  INVX1 _11476_ (
    .A(multiplier_0.op1_15_ ),
    .Y(_05050_)
  );
  INVX1 _11477_ (
    .A(multiplier_0.op2_7_ ),
    .Y(_05051_)
  );
  INVX1 _11478_ (
    .A(multiplier_0.op2_6_ ),
    .Y(_05052_)
  );
  INVX1 _11479_ (
    .A(multiplier_0.op2_5_ ),
    .Y(_05053_)
  );
  INVX1 _11480_ (
    .A(multiplier_0.op2_4_ ),
    .Y(_05054_)
  );
  INVX1 _11481_ (
    .A(multiplier_0.op2_3_ ),
    .Y(_05055_)
  );
  INVX1 _11482_ (
    .A(multiplier_0.op2_2_ ),
    .Y(_05056_)
  );
  INVX1 _11483_ (
    .A(multiplier_0.op2_1_ ),
    .Y(_05057_)
  );
  INVX1 _11484_ (
    .A(multiplier_0.op2_0_ ),
    .Y(_05058_)
  );
  INVX1 _11485_ (
    .A(multiplier_0.op1_6_ ),
    .Y(_05059_)
  );
  INVX1 _11486_ (
    .A(multiplier_0.op1_5_ ),
    .Y(_05060_)
  );
  INVX1 _11487_ (
    .A(multiplier_0.op1_4_ ),
    .Y(_05061_)
  );
  INVX1 _11488_ (
    .A(multiplier_0.op1_3_ ),
    .Y(_05062_)
  );
  INVX1 _11489_ (
    .A(multiplier_0.op1_2_ ),
    .Y(_05063_)
  );
  INVX1 _11490_ (
    .A(multiplier_0.op1_1_ ),
    .Y(_05064_)
  );
  INVX1 _11491_ (
    .A(multiplier_0.op1_0_ ),
    .Y(_05065_)
  );
  INVX1 _11492_ (
    .A(multiplier_0.reshi_13_ ),
    .Y(_05066_)
  );
  INVX1 _11493_ (
    .A(multiplier_0.reshi_11_ ),
    .Y(_05067_)
  );
  INVX1 _11494_ (
    .A(multiplier_0.reshi_9_ ),
    .Y(_05068_)
  );
  INVX1 _11495_ (
    .A(multiplier_0.reshi_7_ ),
    .Y(_05069_)
  );
  INVX1 _11496_ (
    .A(multiplier_0.reshi_0_ ),
    .Y(_05070_)
  );
  INVX1 _11497_ (
    .A(multiplier_0.reslo_12_ ),
    .Y(_05071_)
  );
  INVX1 _11498_ (
    .A(multiplier_0.reslo_5_ ),
    .Y(_05072_)
  );
  INVX1 _11499_ (
    .A(_00110_),
    .Y(_05073_)
  );
  INVX1 _11500_ (
    .A(_00117_),
    .Y(_05074_)
  );
  INVX1 _11501_ (
    .A(_00118_),
    .Y(_05075_)
  );
  INVX1 _11502_ (
    .A(_00119_),
    .Y(_05076_)
  );
  INVX1 _11503_ (
    .A(_00122_),
    .Y(_05077_)
  );
  INVX1 _11504_ (
    .A(_00123_),
    .Y(_05078_)
  );
  INVX1 _11505_ (
    .A(_00162_),
    .Y(_04441_)
  );
  NAND2X1 _11506_ (
    .A(_05042_),
    .B(_00102_),
    .Y(_05079_)
  );
  OR2X1 _11507_ (
    .A(_00101_),
    .B(_05079_),
    .Y(_05080_)
  );
  OR2X1 _11508_ (
    .A(_00099_),
    .B(1'h0),
    .Y(_05081_)
  );
  NAND2X1 _11509_ (
    .A(_05046_),
    .B(_00126_),
    .Y(_05082_)
  );
  NOR2X1 _11510_ (
    .A(_05081_),
    .B(_05082_),
    .Y(_05083_)
  );
  NOR2X1 _11511_ (
    .A(_00108_),
    .B(_05045_),
    .Y(_05084_)
  );
  NOR2X1 _11512_ (
    .A(_00098_),
    .B(_00109_),
    .Y(_05085_)
  );
  NAND2X1 _11513_ (
    .A(_05084_),
    .B(_05085_),
    .Y(_05086_)
  );
  NOR2X1 _11514_ (
    .A(_00106_),
    .B(_00105_),
    .Y(_05087_)
  );
  NAND3X1 _11515_ (
    .A(_00104_),
    .B(_00103_),
    .C(_05087_),
    .Y(_05088_)
  );
  NOR2X1 _11516_ (
    .A(_05086_),
    .B(_05088_),
    .Y(_05089_)
  );
  AND2X1 _11517_ (
    .A(_05083_),
    .B(_05089_),
    .Y(_05090_)
  );
  NOR2X1 _11518_ (
    .A(_00127_),
    .B(_00128_),
    .Y(_05091_)
  );
  OAI21X1 _11519_ (
    .A(_00127_),
    .B(_00128_),
    .C(_05090_),
    .Y(_05092_)
  );
  OR2X1 _11520_ (
    .A(_05080_),
    .B(_05092_),
    .Y(_05093_)
  );
  INVX1 _11521_ (
    .A(_05093_),
    .Y(multiplier_0.op2_wr )
  );
  NOR2X1 _11522_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .Y(_05094_)
  );
  NAND2X1 _11523_ (
    .A(_05047_),
    .B(_05048_),
    .Y(_05095_)
  );
  NAND2X1 _11524_ (
    .A(_05047_),
    .B(multiplier_0.op2_7_ ),
    .Y(_05096_)
  );
  NAND2X1 _11525_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.op2_15_ ),
    .Y(_05097_)
  );
  OAI21X1 _11526_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05051_),
    .C(_05097_),
    .Y(_05098_)
  );
  AND2X1 _11527_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05098_),
    .Y(_05099_)
  );
  OR2X1 _11528_ (
    .A(_05049_),
    .B(_05097_),
    .Y(_05100_)
  );
  NOR2X1 _11529_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05100_),
    .Y(_05101_)
  );
  XNOR2X1 _11530_ (
    .A(_05099_),
    .B(_05101_),
    .Y(_05102_)
  );
  NAND2X1 _11531_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.op2_14_ ),
    .Y(_05103_)
  );
  OAI21X1 _11532_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05052_),
    .C(_05103_),
    .Y(_05104_)
  );
  NAND2X1 _11533_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05104_),
    .Y(_05105_)
  );
  NOR2X1 _11534_ (
    .A(_05102_),
    .B(_05105_),
    .Y(_05106_)
  );
  AOI21X1 _11535_ (
    .A(_05099_),
    .B(_05101_),
    .C(_05106_),
    .Y(_05107_)
  );
  AND2X1 _11536_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05098_),
    .Y(_05108_)
  );
  NOR2X1 _11537_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05100_),
    .Y(_05109_)
  );
  XNOR2X1 _11538_ (
    .A(_05108_),
    .B(_05109_),
    .Y(_05110_)
  );
  NAND2X1 _11539_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05104_),
    .Y(_05111_)
  );
  NOR2X1 _11540_ (
    .A(_05110_),
    .B(_05111_),
    .Y(_05112_)
  );
  XOR2X1 _11541_ (
    .A(_05110_),
    .B(_05111_),
    .Y(_05113_)
  );
  INVX1 _11542_ (
    .A(_05113_),
    .Y(_05114_)
  );
  NOR2X1 _11543_ (
    .A(_05107_),
    .B(_05114_),
    .Y(_05115_)
  );
  XNOR2X1 _11544_ (
    .A(_05107_),
    .B(_05113_),
    .Y(_05116_)
  );
  NAND2X1 _11545_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.op2_11_ ),
    .Y(_05117_)
  );
  OAI21X1 _11546_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05055_),
    .C(_05117_),
    .Y(_05118_)
  );
  NAND2X1 _11547_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05118_),
    .Y(_05119_)
  );
  NAND2X1 _11548_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.op2_12_ ),
    .Y(_05120_)
  );
  MUX2X1 _11549_ (
    .A(multiplier_0.op2_12_ ),
    .B(multiplier_0.op2_4_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05121_)
  );
  OAI21X1 _11550_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05054_),
    .C(_05120_),
    .Y(_05122_)
  );
  NAND2X1 _11551_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05122_),
    .Y(_05123_)
  );
  NAND2X1 _11552_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.op2_13_ ),
    .Y(_05124_)
  );
  MUX2X1 _11553_ (
    .A(multiplier_0.op2_13_ ),
    .B(multiplier_0.op2_5_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05125_)
  );
  OAI21X1 _11554_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05053_),
    .C(_05124_),
    .Y(_05126_)
  );
  NAND2X1 _11555_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05126_),
    .Y(_05127_)
  );
  NAND2X1 _11556_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05126_),
    .Y(_05128_)
  );
  AND2X1 _11557_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05122_),
    .Y(_05129_)
  );
  OR2X1 _11558_ (
    .A(_05123_),
    .B(_05127_),
    .Y(_05130_)
  );
  XNOR2X1 _11559_ (
    .A(_05123_),
    .B(_05127_),
    .Y(_05131_)
  );
  XOR2X1 _11560_ (
    .A(_05119_),
    .B(_05131_),
    .Y(_05132_)
  );
  AOI21X1 _11561_ (
    .A(_05116_),
    .B(_05132_),
    .C(_05115_),
    .Y(_05133_)
  );
  AOI21X1 _11562_ (
    .A(_05108_),
    .B(_05109_),
    .C(_05112_),
    .Y(_05134_)
  );
  AND2X1 _11563_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05098_),
    .Y(_05135_)
  );
  NOR2X1 _11564_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05100_),
    .Y(_05136_)
  );
  XNOR2X1 _11565_ (
    .A(_05135_),
    .B(_05136_),
    .Y(_05137_)
  );
  NAND2X1 _11566_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05104_),
    .Y(_05138_)
  );
  NOR2X1 _11567_ (
    .A(_05137_),
    .B(_05138_),
    .Y(_05139_)
  );
  XOR2X1 _11568_ (
    .A(_05137_),
    .B(_05138_),
    .Y(_05140_)
  );
  INVX1 _11569_ (
    .A(_05140_),
    .Y(_05141_)
  );
  NOR2X1 _11570_ (
    .A(_05134_),
    .B(_05141_),
    .Y(_05142_)
  );
  XNOR2X1 _11571_ (
    .A(_05134_),
    .B(_05140_),
    .Y(_05143_)
  );
  NAND2X1 _11572_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05126_),
    .Y(_05144_)
  );
  OAI21X1 _11573_ (
    .A(_05050_),
    .B(_05121_),
    .C(_05128_),
    .Y(_05145_)
  );
  OAI21X1 _11574_ (
    .A(_05123_),
    .B(_05144_),
    .C(_05145_),
    .Y(_05146_)
  );
  INVX1 _11575_ (
    .A(_05146_),
    .Y(_05147_)
  );
  NOR2X1 _11576_ (
    .A(_05049_),
    .B(_05050_),
    .Y(_05148_)
  );
  NAND2X1 _11577_ (
    .A(multiplier_0.sign_sel ),
    .B(multiplier_0.op1_15_ ),
    .Y(_05149_)
  );
  NOR2X1 _11578_ (
    .A(_05049_),
    .B(_05119_),
    .Y(_05150_)
  );
  NAND2X1 _11579_ (
    .A(_05147_),
    .B(_05150_),
    .Y(_05151_)
  );
  XNOR2X1 _11580_ (
    .A(_05146_),
    .B(_05150_),
    .Y(_05152_)
  );
  AND2X1 _11581_ (
    .A(_05143_),
    .B(_05152_),
    .Y(_05153_)
  );
  XNOR2X1 _11582_ (
    .A(_05143_),
    .B(_05152_),
    .Y(_05154_)
  );
  NOR2X1 _11583_ (
    .A(_05133_),
    .B(_05154_),
    .Y(_05155_)
  );
  XOR2X1 _11584_ (
    .A(_05133_),
    .B(_05154_),
    .Y(_05156_)
  );
  NAND2X1 _11585_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.op2_9_ ),
    .Y(_05157_)
  );
  MUX2X1 _11586_ (
    .A(multiplier_0.op2_9_ ),
    .B(multiplier_0.op2_1_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05158_)
  );
  OAI21X1 _11587_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05057_),
    .C(_05157_),
    .Y(_05159_)
  );
  NOR2X1 _11588_ (
    .A(_05050_),
    .B(_05158_),
    .Y(_05160_)
  );
  NOR2X1 _11589_ (
    .A(_05149_),
    .B(_05158_),
    .Y(_05161_)
  );
  NAND2X1 _11590_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.op2_10_ ),
    .Y(_05162_)
  );
  MUX2X1 _11591_ (
    .A(multiplier_0.op2_10_ ),
    .B(multiplier_0.op2_2_ ),
    .S(multiplier_0.cycle_0_ ),
    .Y(_05163_)
  );
  OAI21X1 _11592_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05056_),
    .C(_05162_),
    .Y(_05164_)
  );
  NOR2X1 _11593_ (
    .A(_05050_),
    .B(_05163_),
    .Y(_05165_)
  );
  NAND2X1 _11594_ (
    .A(_05161_),
    .B(_05164_),
    .Y(_05166_)
  );
  NAND2X1 _11595_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.op2_8_ ),
    .Y(_05167_)
  );
  NAND2X1 _11596_ (
    .A(_05047_),
    .B(multiplier_0.op2_0_ ),
    .Y(_05168_)
  );
  OAI21X1 _11597_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_05058_),
    .C(_05167_),
    .Y(_05169_)
  );
  NAND2X1 _11598_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05169_),
    .Y(_05170_)
  );
  NAND2X1 _11599_ (
    .A(_05148_),
    .B(_05169_),
    .Y(_05171_)
  );
  OAI21X1 _11600_ (
    .A(_05161_),
    .B(_05165_),
    .C(_05166_),
    .Y(_05172_)
  );
  OAI21X1 _11601_ (
    .A(_05171_),
    .B(_05172_),
    .C(_05166_),
    .Y(_05173_)
  );
  INVX1 _11602_ (
    .A(_05173_),
    .Y(_05174_)
  );
  OAI21X1 _11603_ (
    .A(_05119_),
    .B(_05131_),
    .C(_05130_),
    .Y(_05175_)
  );
  NAND3X1 _11604_ (
    .A(_05148_),
    .B(_05169_),
    .C(_05172_),
    .Y(_05176_)
  );
  OAI21X1 _11605_ (
    .A(_05159_),
    .B(_05164_),
    .C(_05148_),
    .Y(_05177_)
  );
  OAI21X1 _11606_ (
    .A(_05173_),
    .B(_05177_),
    .C(_05176_),
    .Y(_05178_)
  );
  XOR2X1 _11607_ (
    .A(_05175_),
    .B(_05178_),
    .Y(_05179_)
  );
  AND2X1 _11608_ (
    .A(_05173_),
    .B(_05179_),
    .Y(_05180_)
  );
  NOR2X1 _11609_ (
    .A(_05173_),
    .B(_05179_),
    .Y(_05181_)
  );
  NOR2X1 _11610_ (
    .A(_05180_),
    .B(_05181_),
    .Y(_05182_)
  );
  AOI21X1 _11611_ (
    .A(_05156_),
    .B(_05182_),
    .C(_05155_),
    .Y(_05183_)
  );
  NOR2X1 _11612_ (
    .A(_05142_),
    .B(_05153_),
    .Y(_05184_)
  );
  AOI21X1 _11613_ (
    .A(_05135_),
    .B(_05136_),
    .C(_05139_),
    .Y(_05185_)
  );
  AND2X1 _11614_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05098_),
    .Y(_05186_)
  );
  NOR2X1 _11615_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05100_),
    .Y(_05187_)
  );
  AND2X1 _11616_ (
    .A(_05186_),
    .B(_05187_),
    .Y(_05188_)
  );
  XNOR2X1 _11617_ (
    .A(_05186_),
    .B(_05187_),
    .Y(_05189_)
  );
  NAND2X1 _11618_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05104_),
    .Y(_05190_)
  );
  NOR2X1 _11619_ (
    .A(_05189_),
    .B(_05190_),
    .Y(_05191_)
  );
  XOR2X1 _11620_ (
    .A(_05189_),
    .B(_05190_),
    .Y(_05192_)
  );
  INVX1 _11621_ (
    .A(_05192_),
    .Y(_05193_)
  );
  NOR2X1 _11622_ (
    .A(_05185_),
    .B(_05193_),
    .Y(_05194_)
  );
  XNOR2X1 _11623_ (
    .A(_05185_),
    .B(_05192_),
    .Y(_05195_)
  );
  OAI21X1 _11624_ (
    .A(_05121_),
    .B(_05149_),
    .C(_05144_),
    .Y(_05196_)
  );
  NAND3X1 _11625_ (
    .A(_05122_),
    .B(_05126_),
    .C(_05148_),
    .Y(_05197_)
  );
  INVX1 _11626_ (
    .A(_05197_),
    .Y(_05198_)
  );
  NAND2X1 _11627_ (
    .A(_05196_),
    .B(_05197_),
    .Y(_05199_)
  );
  NAND2X1 _11628_ (
    .A(_05150_),
    .B(_05199_),
    .Y(_05200_)
  );
  XNOR2X1 _11629_ (
    .A(_05150_),
    .B(_05199_),
    .Y(_05201_)
  );
  AND2X1 _11630_ (
    .A(_05195_),
    .B(_05201_),
    .Y(_05202_)
  );
  NOR2X1 _11631_ (
    .A(_05195_),
    .B(_05201_),
    .Y(_05203_)
  );
  NOR2X1 _11632_ (
    .A(_05202_),
    .B(_05203_),
    .Y(_05204_)
  );
  OAI21X1 _11633_ (
    .A(_05142_),
    .B(_05153_),
    .C(_05204_),
    .Y(_05205_)
  );
  INVX1 _11634_ (
    .A(_05205_),
    .Y(_05206_)
  );
  XNOR2X1 _11635_ (
    .A(_05184_),
    .B(_05204_),
    .Y(_05207_)
  );
  OAI21X1 _11636_ (
    .A(_05123_),
    .B(_05144_),
    .C(_05151_),
    .Y(_05208_)
  );
  AND2X1 _11637_ (
    .A(_05178_),
    .B(_05208_),
    .Y(_05209_)
  );
  NOR2X1 _11638_ (
    .A(_05178_),
    .B(_05208_),
    .Y(_05210_)
  );
  NOR2X1 _11639_ (
    .A(_05209_),
    .B(_05210_),
    .Y(_05211_)
  );
  XNOR2X1 _11640_ (
    .A(_05174_),
    .B(_05211_),
    .Y(_05212_)
  );
  XNOR2X1 _11641_ (
    .A(_05207_),
    .B(_05212_),
    .Y(_05213_)
  );
  NOR2X1 _11642_ (
    .A(_05183_),
    .B(_05213_),
    .Y(_05214_)
  );
  XOR2X1 _11643_ (
    .A(_05183_),
    .B(_05213_),
    .Y(_05215_)
  );
  INVX1 _11644_ (
    .A(_05215_),
    .Y(_05216_)
  );
  AOI21X1 _11645_ (
    .A(_05175_),
    .B(_05178_),
    .C(_05180_),
    .Y(_05217_)
  );
  NOR2X1 _11646_ (
    .A(_05216_),
    .B(_05217_),
    .Y(_05218_)
  );
  NOR2X1 _11647_ (
    .A(_05214_),
    .B(_05218_),
    .Y(_05219_)
  );
  AOI21X1 _11648_ (
    .A(_05207_),
    .B(_05212_),
    .C(_05206_),
    .Y(_05220_)
  );
  NOR2X1 _11649_ (
    .A(_05194_),
    .B(_05202_),
    .Y(_05221_)
  );
  NOR2X1 _11650_ (
    .A(_05188_),
    .B(_05191_),
    .Y(_05222_)
  );
  NAND2X1 _11651_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05098_),
    .Y(_05223_)
  );
  NOR2X1 _11652_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05100_),
    .Y(_05224_)
  );
  NAND3X1 _11653_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05098_),
    .C(_05224_),
    .Y(_05225_)
  );
  OAI21X1 _11654_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05100_),
    .C(_05223_),
    .Y(_05226_)
  );
  NAND2X1 _11655_ (
    .A(_05225_),
    .B(_05226_),
    .Y(_05227_)
  );
  NAND2X1 _11656_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05104_),
    .Y(_05228_)
  );
  OR2X1 _11657_ (
    .A(_05227_),
    .B(_05228_),
    .Y(_05229_)
  );
  XOR2X1 _11658_ (
    .A(_05227_),
    .B(_05228_),
    .Y(_05230_)
  );
  OAI21X1 _11659_ (
    .A(_05188_),
    .B(_05191_),
    .C(_05230_),
    .Y(_05231_)
  );
  XNOR2X1 _11660_ (
    .A(_05222_),
    .B(_05230_),
    .Y(_05232_)
  );
  AOI21X1 _11661_ (
    .A(_05150_),
    .B(_05196_),
    .C(_05198_),
    .Y(_05233_)
  );
  INVX1 _11662_ (
    .A(_05233_),
    .Y(_05234_)
  );
  OAI21X1 _11663_ (
    .A(_05122_),
    .B(_05126_),
    .C(_05148_),
    .Y(_05235_)
  );
  OAI21X1 _11664_ (
    .A(_05234_),
    .B(_05235_),
    .C(_05200_),
    .Y(_05236_)
  );
  NAND2X1 _11665_ (
    .A(_05232_),
    .B(_05236_),
    .Y(_05237_)
  );
  XOR2X1 _11666_ (
    .A(_05232_),
    .B(_05236_),
    .Y(_05238_)
  );
  OAI21X1 _11667_ (
    .A(_05194_),
    .B(_05202_),
    .C(_05238_),
    .Y(_05239_)
  );
  XNOR2X1 _11668_ (
    .A(_05221_),
    .B(_05238_),
    .Y(_05240_)
  );
  XNOR2X1 _11669_ (
    .A(_05178_),
    .B(_05234_),
    .Y(_05241_)
  );
  NOR2X1 _11670_ (
    .A(_05174_),
    .B(_05241_),
    .Y(_05242_)
  );
  XNOR2X1 _11671_ (
    .A(_05173_),
    .B(_05241_),
    .Y(_05243_)
  );
  NAND2X1 _11672_ (
    .A(_05240_),
    .B(_05243_),
    .Y(_05244_)
  );
  XNOR2X1 _11673_ (
    .A(_05240_),
    .B(_05243_),
    .Y(_05245_)
  );
  NOR2X1 _11674_ (
    .A(_05220_),
    .B(_05245_),
    .Y(_05246_)
  );
  XOR2X1 _11675_ (
    .A(_05220_),
    .B(_05245_),
    .Y(_05247_)
  );
  INVX1 _11676_ (
    .A(_05247_),
    .Y(_05248_)
  );
  AOI21X1 _11677_ (
    .A(_05173_),
    .B(_05211_),
    .C(_05209_),
    .Y(_05249_)
  );
  NOR2X1 _11678_ (
    .A(_05248_),
    .B(_05249_),
    .Y(_05250_)
  );
  XNOR2X1 _11679_ (
    .A(_05247_),
    .B(_05249_),
    .Y(_05251_)
  );
  OAI21X1 _11680_ (
    .A(_05214_),
    .B(_05218_),
    .C(_05251_),
    .Y(_05252_)
  );
  NOR2X1 _11681_ (
    .A(_05246_),
    .B(_05250_),
    .Y(_05253_)
  );
  NAND2X1 _11682_ (
    .A(_05231_),
    .B(_05237_),
    .Y(_05254_)
  );
  NAND2X1 _11683_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05098_),
    .Y(_05255_)
  );
  NOR2X1 _11684_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05100_),
    .Y(_05256_)
  );
  OAI21X1 _11685_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05100_),
    .C(_05255_),
    .Y(_05257_)
  );
  NAND3X1 _11686_ (
    .A(multiplier_0.op1_15_ ),
    .B(_05098_),
    .C(_05256_),
    .Y(_05258_)
  );
  NAND2X1 _11687_ (
    .A(_05257_),
    .B(_05258_),
    .Y(_05259_)
  );
  NAND2X1 _11688_ (
    .A(_05104_),
    .B(_05148_),
    .Y(_05260_)
  );
  XNOR2X1 _11689_ (
    .A(_05259_),
    .B(_05260_),
    .Y(_05261_)
  );
  AOI21X1 _11690_ (
    .A(_05225_),
    .B(_05229_),
    .C(_05261_),
    .Y(_05262_)
  );
  INVX1 _11691_ (
    .A(_05262_),
    .Y(_05263_)
  );
  NAND3X1 _11692_ (
    .A(_05225_),
    .B(_05229_),
    .C(_05261_),
    .Y(_05264_)
  );
  AND2X1 _11693_ (
    .A(_05263_),
    .B(_05264_),
    .Y(_05265_)
  );
  XNOR2X1 _11694_ (
    .A(_05236_),
    .B(_05265_),
    .Y(_05266_)
  );
  AOI21X1 _11695_ (
    .A(_05231_),
    .B(_05237_),
    .C(_05266_),
    .Y(_05267_)
  );
  XOR2X1 _11696_ (
    .A(_05254_),
    .B(_05266_),
    .Y(_05268_)
  );
  INVX1 _11697_ (
    .A(_05268_),
    .Y(_05269_)
  );
  XOR2X1 _11698_ (
    .A(_05243_),
    .B(_05268_),
    .Y(_05270_)
  );
  NAND3X1 _11699_ (
    .A(_05239_),
    .B(_05244_),
    .C(_05270_),
    .Y(_05271_)
  );
  AOI21X1 _11700_ (
    .A(_05239_),
    .B(_05244_),
    .C(_05270_),
    .Y(_05272_)
  );
  INVX1 _11701_ (
    .A(_05272_),
    .Y(_05273_)
  );
  NAND2X1 _11702_ (
    .A(_05271_),
    .B(_05273_),
    .Y(_05274_)
  );
  AOI21X1 _11703_ (
    .A(_05178_),
    .B(_05234_),
    .C(_05242_),
    .Y(_05275_)
  );
  XNOR2X1 _11704_ (
    .A(_05274_),
    .B(_05275_),
    .Y(_05276_)
  );
  NOR2X1 _11705_ (
    .A(_05253_),
    .B(_05276_),
    .Y(_05277_)
  );
  XNOR2X1 _11706_ (
    .A(_05253_),
    .B(_05276_),
    .Y(_05278_)
  );
  NOR2X1 _11707_ (
    .A(_05252_),
    .B(_05278_),
    .Y(_05279_)
  );
  AND2X1 _11708_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05098_),
    .Y(_05280_)
  );
  NOR2X1 _11709_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05100_),
    .Y(_05281_)
  );
  XNOR2X1 _11710_ (
    .A(_05280_),
    .B(_05281_),
    .Y(_05282_)
  );
  NAND2X1 _11711_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05104_),
    .Y(_05283_)
  );
  NOR2X1 _11712_ (
    .A(_05282_),
    .B(_05283_),
    .Y(_05284_)
  );
  AOI21X1 _11713_ (
    .A(_05280_),
    .B(_05281_),
    .C(_05284_),
    .Y(_05285_)
  );
  XOR2X1 _11714_ (
    .A(_05102_),
    .B(_05105_),
    .Y(_05286_)
  );
  INVX1 _11715_ (
    .A(_05286_),
    .Y(_05287_)
  );
  NOR2X1 _11716_ (
    .A(_05285_),
    .B(_05287_),
    .Y(_05288_)
  );
  XNOR2X1 _11717_ (
    .A(_05285_),
    .B(_05286_),
    .Y(_05289_)
  );
  NAND2X1 _11718_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05118_),
    .Y(_05290_)
  );
  NAND2X1 _11719_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05126_),
    .Y(_05291_)
  );
  AND2X1 _11720_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05122_),
    .Y(_05292_)
  );
  NAND3X1 _11721_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05126_),
    .C(_05129_),
    .Y(_05293_)
  );
  XOR2X1 _11722_ (
    .A(_05129_),
    .B(_05291_),
    .Y(_05294_)
  );
  XOR2X1 _11723_ (
    .A(_05290_),
    .B(_05294_),
    .Y(_05295_)
  );
  AOI21X1 _11724_ (
    .A(_05289_),
    .B(_05295_),
    .C(_05288_),
    .Y(_05296_)
  );
  XNOR2X1 _11725_ (
    .A(_05116_),
    .B(_05132_),
    .Y(_05297_)
  );
  NOR2X1 _11726_ (
    .A(_05296_),
    .B(_05297_),
    .Y(_05298_)
  );
  XOR2X1 _11727_ (
    .A(_05296_),
    .B(_05297_),
    .Y(_05299_)
  );
  OAI21X1 _11728_ (
    .A(_05290_),
    .B(_05294_),
    .C(_05293_),
    .Y(_05300_)
  );
  XOR2X1 _11729_ (
    .A(_05178_),
    .B(_05300_),
    .Y(_05301_)
  );
  AND2X1 _11730_ (
    .A(_05173_),
    .B(_05301_),
    .Y(_05302_)
  );
  NOR2X1 _11731_ (
    .A(_05173_),
    .B(_05301_),
    .Y(_05303_)
  );
  NOR2X1 _11732_ (
    .A(_05302_),
    .B(_05303_),
    .Y(_05304_)
  );
  AOI21X1 _11733_ (
    .A(_05299_),
    .B(_05304_),
    .C(_05298_),
    .Y(_05305_)
  );
  XNOR2X1 _11734_ (
    .A(_05156_),
    .B(_05182_),
    .Y(_05306_)
  );
  NOR2X1 _11735_ (
    .A(_05305_),
    .B(_05306_),
    .Y(_05307_)
  );
  XOR2X1 _11736_ (
    .A(_05305_),
    .B(_05306_),
    .Y(_05308_)
  );
  AOI21X1 _11737_ (
    .A(_05178_),
    .B(_05300_),
    .C(_05302_),
    .Y(_05309_)
  );
  INVX1 _11738_ (
    .A(_05309_),
    .Y(_05310_)
  );
  AOI21X1 _11739_ (
    .A(_05308_),
    .B(_05310_),
    .C(_05307_),
    .Y(_05311_)
  );
  INVX1 _11740_ (
    .A(_05311_),
    .Y(_05312_)
  );
  XNOR2X1 _11741_ (
    .A(_05215_),
    .B(_05217_),
    .Y(_05313_)
  );
  NAND2X1 _11742_ (
    .A(_05312_),
    .B(_05313_),
    .Y(_05314_)
  );
  XNOR2X1 _11743_ (
    .A(_05219_),
    .B(_05251_),
    .Y(_05315_)
  );
  NAND3X1 _11744_ (
    .A(_05312_),
    .B(_05313_),
    .C(_05315_),
    .Y(_05316_)
  );
  AND2X1 _11745_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05098_),
    .Y(_05317_)
  );
  NOR2X1 _11746_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05100_),
    .Y(_05318_)
  );
  XNOR2X1 _11747_ (
    .A(_05317_),
    .B(_05318_),
    .Y(_05319_)
  );
  NAND2X1 _11748_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05104_),
    .Y(_05320_)
  );
  NOR2X1 _11749_ (
    .A(_05319_),
    .B(_05320_),
    .Y(_05321_)
  );
  AOI21X1 _11750_ (
    .A(_05317_),
    .B(_05318_),
    .C(_05321_),
    .Y(_05322_)
  );
  XOR2X1 _11751_ (
    .A(_05282_),
    .B(_05283_),
    .Y(_05323_)
  );
  INVX1 _11752_ (
    .A(_05323_),
    .Y(_05324_)
  );
  NOR2X1 _11753_ (
    .A(_05322_),
    .B(_05324_),
    .Y(_05325_)
  );
  XNOR2X1 _11754_ (
    .A(_05322_),
    .B(_05323_),
    .Y(_05326_)
  );
  NAND2X1 _11755_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05118_),
    .Y(_05327_)
  );
  NAND2X1 _11756_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05126_),
    .Y(_05328_)
  );
  AND2X1 _11757_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05122_),
    .Y(_05329_)
  );
  NAND3X1 _11758_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05126_),
    .C(_05292_),
    .Y(_05330_)
  );
  XOR2X1 _11759_ (
    .A(_05292_),
    .B(_05328_),
    .Y(_05331_)
  );
  XOR2X1 _11760_ (
    .A(_05327_),
    .B(_05331_),
    .Y(_05332_)
  );
  AOI21X1 _11761_ (
    .A(_05326_),
    .B(_05332_),
    .C(_05325_),
    .Y(_05333_)
  );
  XNOR2X1 _11762_ (
    .A(_05289_),
    .B(_05295_),
    .Y(_05334_)
  );
  OR2X1 _11763_ (
    .A(_05333_),
    .B(_05334_),
    .Y(_05335_)
  );
  NAND2X1 _11764_ (
    .A(_05333_),
    .B(_05334_),
    .Y(_05336_)
  );
  NAND2X1 _11765_ (
    .A(_05335_),
    .B(_05336_),
    .Y(_05337_)
  );
  NAND2X1 _11766_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05164_),
    .Y(_05338_)
  );
  AND2X1 _11767_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05159_),
    .Y(_05339_)
  );
  NAND3X1 _11768_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05160_),
    .C(_05164_),
    .Y(_05340_)
  );
  XOR2X1 _11769_ (
    .A(_05160_),
    .B(_05338_),
    .Y(_05341_)
  );
  OAI21X1 _11770_ (
    .A(_05171_),
    .B(_05341_),
    .C(_05340_),
    .Y(_05342_)
  );
  OAI21X1 _11771_ (
    .A(_05327_),
    .B(_05331_),
    .C(_05330_),
    .Y(_05343_)
  );
  INVX1 _11772_ (
    .A(_05343_),
    .Y(_05344_)
  );
  XNOR2X1 _11773_ (
    .A(_05171_),
    .B(_05172_),
    .Y(_05345_)
  );
  XNOR2X1 _11774_ (
    .A(_05343_),
    .B(_05345_),
    .Y(_05346_)
  );
  NAND2X1 _11775_ (
    .A(_05342_),
    .B(_05346_),
    .Y(_05347_)
  );
  XNOR2X1 _11776_ (
    .A(_05342_),
    .B(_05346_),
    .Y(_05348_)
  );
  OAI21X1 _11777_ (
    .A(_05337_),
    .B(_05348_),
    .C(_05335_),
    .Y(_05349_)
  );
  INVX1 _11778_ (
    .A(_05349_),
    .Y(_05350_)
  );
  XNOR2X1 _11779_ (
    .A(_05299_),
    .B(_05304_),
    .Y(_05351_)
  );
  NOR2X1 _11780_ (
    .A(_05350_),
    .B(_05351_),
    .Y(_05352_)
  );
  OAI21X1 _11781_ (
    .A(_05344_),
    .B(_05345_),
    .C(_05347_),
    .Y(_05353_)
  );
  INVX1 _11782_ (
    .A(_05353_),
    .Y(_05354_)
  );
  XOR2X1 _11783_ (
    .A(_05349_),
    .B(_05351_),
    .Y(_05355_)
  );
  NOR2X1 _11784_ (
    .A(_05354_),
    .B(_05355_),
    .Y(_05356_)
  );
  NOR2X1 _11785_ (
    .A(_05352_),
    .B(_05356_),
    .Y(_05357_)
  );
  XNOR2X1 _11786_ (
    .A(_05308_),
    .B(_05309_),
    .Y(_05358_)
  );
  OAI21X1 _11787_ (
    .A(_05352_),
    .B(_05356_),
    .C(_05358_),
    .Y(_05359_)
  );
  XNOR2X1 _11788_ (
    .A(_05312_),
    .B(_05313_),
    .Y(_05360_)
  );
  NOR2X1 _11789_ (
    .A(_05359_),
    .B(_05360_),
    .Y(_05361_)
  );
  AND2X1 _11790_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05098_),
    .Y(_05362_)
  );
  NOR2X1 _11791_ (
    .A(multiplier_0.op1_6_ ),
    .B(_05100_),
    .Y(_05363_)
  );
  NAND2X1 _11792_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05104_),
    .Y(_05364_)
  );
  XNOR2X1 _11793_ (
    .A(_05362_),
    .B(_05363_),
    .Y(_05365_)
  );
  NOR2X1 _11794_ (
    .A(_05364_),
    .B(_05365_),
    .Y(_05366_)
  );
  AOI21X1 _11795_ (
    .A(_05362_),
    .B(_05363_),
    .C(_05366_),
    .Y(_05367_)
  );
  XOR2X1 _11796_ (
    .A(_05319_),
    .B(_05320_),
    .Y(_05368_)
  );
  INVX1 _11797_ (
    .A(_05368_),
    .Y(_05369_)
  );
  NOR2X1 _11798_ (
    .A(_05367_),
    .B(_05369_),
    .Y(_05370_)
  );
  XNOR2X1 _11799_ (
    .A(_05367_),
    .B(_05368_),
    .Y(_05371_)
  );
  NAND2X1 _11800_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05118_),
    .Y(_05372_)
  );
  NAND2X1 _11801_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05126_),
    .Y(_05373_)
  );
  AND2X1 _11802_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05122_),
    .Y(_05374_)
  );
  NAND3X1 _11803_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05126_),
    .C(_05329_),
    .Y(_05375_)
  );
  XOR2X1 _11804_ (
    .A(_05329_),
    .B(_05373_),
    .Y(_05376_)
  );
  XOR2X1 _11805_ (
    .A(_05372_),
    .B(_05376_),
    .Y(_05377_)
  );
  AOI21X1 _11806_ (
    .A(_05371_),
    .B(_05377_),
    .C(_05370_),
    .Y(_05378_)
  );
  XNOR2X1 _11807_ (
    .A(_05326_),
    .B(_05332_),
    .Y(_05379_)
  );
  OR2X1 _11808_ (
    .A(_05378_),
    .B(_05379_),
    .Y(_05380_)
  );
  NAND2X1 _11809_ (
    .A(_05378_),
    .B(_05379_),
    .Y(_05381_)
  );
  NAND2X1 _11810_ (
    .A(_05380_),
    .B(_05381_),
    .Y(_05382_)
  );
  NAND2X1 _11811_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05164_),
    .Y(_05383_)
  );
  AND2X1 _11812_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05159_),
    .Y(_05384_)
  );
  NAND3X1 _11813_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05164_),
    .C(_05339_),
    .Y(_05385_)
  );
  XOR2X1 _11814_ (
    .A(_05339_),
    .B(_05383_),
    .Y(_05386_)
  );
  OAI21X1 _11815_ (
    .A(_05170_),
    .B(_05386_),
    .C(_05385_),
    .Y(_05387_)
  );
  XNOR2X1 _11816_ (
    .A(_05171_),
    .B(_05341_),
    .Y(_05388_)
  );
  INVX1 _11817_ (
    .A(_05388_),
    .Y(_05389_)
  );
  OAI21X1 _11818_ (
    .A(_05372_),
    .B(_05376_),
    .C(_05375_),
    .Y(_05390_)
  );
  NAND2X1 _11819_ (
    .A(_05389_),
    .B(_05390_),
    .Y(_05391_)
  );
  XOR2X1 _11820_ (
    .A(_05388_),
    .B(_05390_),
    .Y(_05392_)
  );
  INVX1 _11821_ (
    .A(_05392_),
    .Y(_05393_)
  );
  NAND2X1 _11822_ (
    .A(_05387_),
    .B(_05393_),
    .Y(_05394_)
  );
  XOR2X1 _11823_ (
    .A(_05387_),
    .B(_05392_),
    .Y(_05395_)
  );
  OAI21X1 _11824_ (
    .A(_05382_),
    .B(_05395_),
    .C(_05380_),
    .Y(_05396_)
  );
  INVX1 _11825_ (
    .A(_05396_),
    .Y(_05397_)
  );
  XNOR2X1 _11826_ (
    .A(_05337_),
    .B(_05348_),
    .Y(_05398_)
  );
  XOR2X1 _11827_ (
    .A(_05396_),
    .B(_05398_),
    .Y(_05399_)
  );
  AOI21X1 _11828_ (
    .A(_05391_),
    .B(_05394_),
    .C(_05399_),
    .Y(_05400_)
  );
  INVX1 _11829_ (
    .A(_05400_),
    .Y(_05401_)
  );
  OAI21X1 _11830_ (
    .A(_05397_),
    .B(_05398_),
    .C(_05401_),
    .Y(_05402_)
  );
  XNOR2X1 _11831_ (
    .A(_05354_),
    .B(_05355_),
    .Y(_05403_)
  );
  INVX1 _11832_ (
    .A(_05403_),
    .Y(_05404_)
  );
  NAND2X1 _11833_ (
    .A(_05402_),
    .B(_05404_),
    .Y(_05405_)
  );
  XOR2X1 _11834_ (
    .A(_05357_),
    .B(_05358_),
    .Y(_05406_)
  );
  OR2X1 _11835_ (
    .A(_05405_),
    .B(_05406_),
    .Y(_05407_)
  );
  XOR2X1 _11836_ (
    .A(_05405_),
    .B(_05406_),
    .Y(_05408_)
  );
  INVX1 _11837_ (
    .A(_05408_),
    .Y(_05409_)
  );
  AND2X1 _11838_ (
    .A(multiplier_0.op1_6_ ),
    .B(_05098_),
    .Y(_05410_)
  );
  NOR2X1 _11839_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05100_),
    .Y(_05411_)
  );
  NAND2X1 _11840_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05104_),
    .Y(_05412_)
  );
  XNOR2X1 _11841_ (
    .A(_05410_),
    .B(_05411_),
    .Y(_05413_)
  );
  NOR2X1 _11842_ (
    .A(_05412_),
    .B(_05413_),
    .Y(_05414_)
  );
  AOI21X1 _11843_ (
    .A(_05410_),
    .B(_05411_),
    .C(_05414_),
    .Y(_05415_)
  );
  XNOR2X1 _11844_ (
    .A(_05364_),
    .B(_05365_),
    .Y(_05416_)
  );
  NOR2X1 _11845_ (
    .A(_05415_),
    .B(_05416_),
    .Y(_05417_)
  );
  XOR2X1 _11846_ (
    .A(_05415_),
    .B(_05416_),
    .Y(_05418_)
  );
  NAND2X1 _11847_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05118_),
    .Y(_05419_)
  );
  NAND2X1 _11848_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05126_),
    .Y(_05420_)
  );
  AND2X1 _11849_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05122_),
    .Y(_05421_)
  );
  NAND3X1 _11850_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05126_),
    .C(_05374_),
    .Y(_05422_)
  );
  XOR2X1 _11851_ (
    .A(_05374_),
    .B(_05420_),
    .Y(_05423_)
  );
  XOR2X1 _11852_ (
    .A(_05419_),
    .B(_05423_),
    .Y(_05424_)
  );
  AOI21X1 _11853_ (
    .A(_05418_),
    .B(_05424_),
    .C(_05417_),
    .Y(_05425_)
  );
  XNOR2X1 _11854_ (
    .A(_05371_),
    .B(_05377_),
    .Y(_05426_)
  );
  NOR2X1 _11855_ (
    .A(_05425_),
    .B(_05426_),
    .Y(_05427_)
  );
  XOR2X1 _11856_ (
    .A(_05425_),
    .B(_05426_),
    .Y(_05428_)
  );
  NAND2X1 _11857_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05164_),
    .Y(_05429_)
  );
  AND2X1 _11858_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05159_),
    .Y(_05430_)
  );
  NAND3X1 _11859_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05164_),
    .C(_05384_),
    .Y(_05431_)
  );
  XOR2X1 _11860_ (
    .A(_05384_),
    .B(_05429_),
    .Y(_05432_)
  );
  NAND2X1 _11861_ (
    .A(multiplier_0.op1_14_ ),
    .B(_05169_),
    .Y(_05433_)
  );
  OAI21X1 _11862_ (
    .A(_05432_),
    .B(_05433_),
    .C(_05431_),
    .Y(_05434_)
  );
  XNOR2X1 _11863_ (
    .A(_05170_),
    .B(_05386_),
    .Y(_05435_)
  );
  OAI21X1 _11864_ (
    .A(_05419_),
    .B(_05423_),
    .C(_05422_),
    .Y(_05436_)
  );
  INVX1 _11865_ (
    .A(_05436_),
    .Y(_05437_)
  );
  XOR2X1 _11866_ (
    .A(_05435_),
    .B(_05436_),
    .Y(_05438_)
  );
  INVX1 _11867_ (
    .A(_05438_),
    .Y(_05439_)
  );
  NAND2X1 _11868_ (
    .A(_05434_),
    .B(_05439_),
    .Y(_05440_)
  );
  XNOR2X1 _11869_ (
    .A(_05434_),
    .B(_05438_),
    .Y(_05441_)
  );
  AOI21X1 _11870_ (
    .A(_05428_),
    .B(_05441_),
    .C(_05427_),
    .Y(_05442_)
  );
  XNOR2X1 _11871_ (
    .A(_05382_),
    .B(_05395_),
    .Y(_05443_)
  );
  OR2X1 _11872_ (
    .A(_05442_),
    .B(_05443_),
    .Y(_05444_)
  );
  XOR2X1 _11873_ (
    .A(_05442_),
    .B(_05443_),
    .Y(_05445_)
  );
  OAI21X1 _11874_ (
    .A(_05435_),
    .B(_05437_),
    .C(_05440_),
    .Y(_05446_)
  );
  NAND2X1 _11875_ (
    .A(_05445_),
    .B(_05446_),
    .Y(_05447_)
  );
  NAND3X1 _11876_ (
    .A(_05391_),
    .B(_05394_),
    .C(_05399_),
    .Y(_05448_)
  );
  NAND2X1 _11877_ (
    .A(_05401_),
    .B(_05448_),
    .Y(_05449_)
  );
  AOI21X1 _11878_ (
    .A(_05444_),
    .B(_05447_),
    .C(_05449_),
    .Y(_05450_)
  );
  INVX1 _11879_ (
    .A(_05450_),
    .Y(_05451_)
  );
  XNOR2X1 _11880_ (
    .A(_05402_),
    .B(_05404_),
    .Y(_05452_)
  );
  NOR2X1 _11881_ (
    .A(_05451_),
    .B(_05452_),
    .Y(_05453_)
  );
  XNOR2X1 _11882_ (
    .A(_05450_),
    .B(_05452_),
    .Y(_05454_)
  );
  AND2X1 _11883_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05098_),
    .Y(_05455_)
  );
  NOR2X1 _11884_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05100_),
    .Y(_05456_)
  );
  NAND2X1 _11885_ (
    .A(multiplier_0.op1_6_ ),
    .B(_05104_),
    .Y(_05457_)
  );
  XNOR2X1 _11886_ (
    .A(_05455_),
    .B(_05456_),
    .Y(_05458_)
  );
  NOR2X1 _11887_ (
    .A(_05457_),
    .B(_05458_),
    .Y(_05459_)
  );
  AOI21X1 _11888_ (
    .A(_05455_),
    .B(_05456_),
    .C(_05459_),
    .Y(_05460_)
  );
  XNOR2X1 _11889_ (
    .A(_05412_),
    .B(_05413_),
    .Y(_05461_)
  );
  NOR2X1 _11890_ (
    .A(_05460_),
    .B(_05461_),
    .Y(_05462_)
  );
  XOR2X1 _11891_ (
    .A(_05460_),
    .B(_05461_),
    .Y(_05463_)
  );
  NAND2X1 _11892_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05118_),
    .Y(_05464_)
  );
  NAND2X1 _11893_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05126_),
    .Y(_05465_)
  );
  AND2X1 _11894_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05122_),
    .Y(_05466_)
  );
  NAND3X1 _11895_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05126_),
    .C(_05421_),
    .Y(_05467_)
  );
  XOR2X1 _11896_ (
    .A(_05421_),
    .B(_05465_),
    .Y(_05468_)
  );
  XOR2X1 _11897_ (
    .A(_05464_),
    .B(_05468_),
    .Y(_05469_)
  );
  AOI21X1 _11898_ (
    .A(_05463_),
    .B(_05469_),
    .C(_05462_),
    .Y(_05470_)
  );
  XNOR2X1 _11899_ (
    .A(_05418_),
    .B(_05424_),
    .Y(_05471_)
  );
  NOR2X1 _11900_ (
    .A(_05470_),
    .B(_05471_),
    .Y(_05472_)
  );
  XOR2X1 _11901_ (
    .A(_05470_),
    .B(_05471_),
    .Y(_05473_)
  );
  NAND2X1 _11902_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05164_),
    .Y(_05474_)
  );
  AND2X1 _11903_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05159_),
    .Y(_05475_)
  );
  NAND3X1 _11904_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05164_),
    .C(_05430_),
    .Y(_05476_)
  );
  XOR2X1 _11905_ (
    .A(_05430_),
    .B(_05474_),
    .Y(_05477_)
  );
  NAND2X1 _11906_ (
    .A(multiplier_0.op1_13_ ),
    .B(_05169_),
    .Y(_05478_)
  );
  OAI21X1 _11907_ (
    .A(_05477_),
    .B(_05478_),
    .C(_05476_),
    .Y(_05479_)
  );
  XOR2X1 _11908_ (
    .A(_05432_),
    .B(_05433_),
    .Y(_05480_)
  );
  OAI21X1 _11909_ (
    .A(_05464_),
    .B(_05468_),
    .C(_05467_),
    .Y(_05481_)
  );
  NAND2X1 _11910_ (
    .A(_05480_),
    .B(_05481_),
    .Y(_05482_)
  );
  XOR2X1 _11911_ (
    .A(_05480_),
    .B(_05481_),
    .Y(_05483_)
  );
  NAND2X1 _11912_ (
    .A(_05479_),
    .B(_05483_),
    .Y(_05484_)
  );
  XOR2X1 _11913_ (
    .A(_05479_),
    .B(_05483_),
    .Y(_05485_)
  );
  AOI21X1 _11914_ (
    .A(_05473_),
    .B(_05485_),
    .C(_05472_),
    .Y(_05486_)
  );
  XNOR2X1 _11915_ (
    .A(_05428_),
    .B(_05441_),
    .Y(_05487_)
  );
  XOR2X1 _11916_ (
    .A(_05486_),
    .B(_05487_),
    .Y(_05488_)
  );
  NAND2X1 _11917_ (
    .A(_05482_),
    .B(_05484_),
    .Y(_05489_)
  );
  NAND2X1 _11918_ (
    .A(_05488_),
    .B(_05489_),
    .Y(_05490_)
  );
  OAI21X1 _11919_ (
    .A(_05486_),
    .B(_05487_),
    .C(_05490_),
    .Y(_05491_)
  );
  XOR2X1 _11920_ (
    .A(_05445_),
    .B(_05446_),
    .Y(_05492_)
  );
  AND2X1 _11921_ (
    .A(_05491_),
    .B(_05492_),
    .Y(_05493_)
  );
  NAND3X1 _11922_ (
    .A(_05444_),
    .B(_05447_),
    .C(_05449_),
    .Y(_05494_)
  );
  AND2X1 _11923_ (
    .A(_05451_),
    .B(_05494_),
    .Y(_05495_)
  );
  NAND2X1 _11924_ (
    .A(_05493_),
    .B(_05495_),
    .Y(_05496_)
  );
  AND2X1 _11925_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05098_),
    .Y(_05497_)
  );
  NOR2X1 _11926_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05100_),
    .Y(_05498_)
  );
  NAND2X1 _11927_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05104_),
    .Y(_05499_)
  );
  XNOR2X1 _11928_ (
    .A(_05497_),
    .B(_05498_),
    .Y(_05500_)
  );
  NOR2X1 _11929_ (
    .A(_05499_),
    .B(_05500_),
    .Y(_05501_)
  );
  AOI21X1 _11930_ (
    .A(_05497_),
    .B(_05498_),
    .C(_05501_),
    .Y(_05502_)
  );
  XNOR2X1 _11931_ (
    .A(_05457_),
    .B(_05458_),
    .Y(_05503_)
  );
  NOR2X1 _11932_ (
    .A(_05502_),
    .B(_05503_),
    .Y(_05504_)
  );
  XOR2X1 _11933_ (
    .A(_05502_),
    .B(_05503_),
    .Y(_05505_)
  );
  NAND2X1 _11934_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05118_),
    .Y(_05506_)
  );
  NAND2X1 _11935_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05126_),
    .Y(_05507_)
  );
  AND2X1 _11936_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05122_),
    .Y(_05508_)
  );
  NAND3X1 _11937_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05126_),
    .C(_05466_),
    .Y(_05509_)
  );
  XOR2X1 _11938_ (
    .A(_05466_),
    .B(_05507_),
    .Y(_05510_)
  );
  XOR2X1 _11939_ (
    .A(_05506_),
    .B(_05510_),
    .Y(_05511_)
  );
  AOI21X1 _11940_ (
    .A(_05505_),
    .B(_05511_),
    .C(_05504_),
    .Y(_05512_)
  );
  XNOR2X1 _11941_ (
    .A(_05463_),
    .B(_05469_),
    .Y(_05513_)
  );
  NOR2X1 _11942_ (
    .A(_05512_),
    .B(_05513_),
    .Y(_05514_)
  );
  XOR2X1 _11943_ (
    .A(_05512_),
    .B(_05513_),
    .Y(_05515_)
  );
  NAND2X1 _11944_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05164_),
    .Y(_05516_)
  );
  AND2X1 _11945_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05159_),
    .Y(_05517_)
  );
  NAND3X1 _11946_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05164_),
    .C(_05475_),
    .Y(_05518_)
  );
  XOR2X1 _11947_ (
    .A(_05475_),
    .B(_05516_),
    .Y(_05519_)
  );
  NAND2X1 _11948_ (
    .A(multiplier_0.op1_12_ ),
    .B(_05169_),
    .Y(_05520_)
  );
  OAI21X1 _11949_ (
    .A(_05519_),
    .B(_05520_),
    .C(_05518_),
    .Y(_05521_)
  );
  XOR2X1 _11950_ (
    .A(_05477_),
    .B(_05478_),
    .Y(_05522_)
  );
  OAI21X1 _11951_ (
    .A(_05506_),
    .B(_05510_),
    .C(_05509_),
    .Y(_05523_)
  );
  NAND2X1 _11952_ (
    .A(_05522_),
    .B(_05523_),
    .Y(_05524_)
  );
  XOR2X1 _11953_ (
    .A(_05522_),
    .B(_05523_),
    .Y(_05525_)
  );
  NAND2X1 _11954_ (
    .A(_05521_),
    .B(_05525_),
    .Y(_05526_)
  );
  XOR2X1 _11955_ (
    .A(_05521_),
    .B(_05525_),
    .Y(_05527_)
  );
  AOI21X1 _11956_ (
    .A(_05515_),
    .B(_05527_),
    .C(_05514_),
    .Y(_05528_)
  );
  XNOR2X1 _11957_ (
    .A(_05473_),
    .B(_05485_),
    .Y(_05529_)
  );
  OR2X1 _11958_ (
    .A(_05528_),
    .B(_05529_),
    .Y(_05530_)
  );
  NAND2X1 _11959_ (
    .A(_05524_),
    .B(_05526_),
    .Y(_05531_)
  );
  XOR2X1 _11960_ (
    .A(_05528_),
    .B(_05529_),
    .Y(_05532_)
  );
  NAND2X1 _11961_ (
    .A(_05531_),
    .B(_05532_),
    .Y(_05533_)
  );
  OAI21X1 _11962_ (
    .A(_05528_),
    .B(_05529_),
    .C(_05533_),
    .Y(_05534_)
  );
  XNOR2X1 _11963_ (
    .A(_05488_),
    .B(_05489_),
    .Y(_05535_)
  );
  AOI21X1 _11964_ (
    .A(_05530_),
    .B(_05533_),
    .C(_05535_),
    .Y(_05536_)
  );
  NOR2X1 _11965_ (
    .A(_05491_),
    .B(_05492_),
    .Y(_05537_)
  );
  NOR2X1 _11966_ (
    .A(_05493_),
    .B(_05537_),
    .Y(_05538_)
  );
  AND2X1 _11967_ (
    .A(_05536_),
    .B(_05538_),
    .Y(_05539_)
  );
  XNOR2X1 _11968_ (
    .A(_05536_),
    .B(_05538_),
    .Y(_05540_)
  );
  INVX1 _11969_ (
    .A(_05540_),
    .Y(_05541_)
  );
  AND2X1 _11970_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05098_),
    .Y(_05542_)
  );
  NOR2X1 _11971_ (
    .A(multiplier_0.op1_2_ ),
    .B(_05100_),
    .Y(_05543_)
  );
  NAND2X1 _11972_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05104_),
    .Y(_05544_)
  );
  XNOR2X1 _11973_ (
    .A(_05542_),
    .B(_05543_),
    .Y(_05545_)
  );
  NOR2X1 _11974_ (
    .A(_05544_),
    .B(_05545_),
    .Y(_05546_)
  );
  AOI21X1 _11975_ (
    .A(_05542_),
    .B(_05543_),
    .C(_05546_),
    .Y(_05547_)
  );
  XNOR2X1 _11976_ (
    .A(_05499_),
    .B(_05500_),
    .Y(_05548_)
  );
  NOR2X1 _11977_ (
    .A(_05547_),
    .B(_05548_),
    .Y(_05549_)
  );
  XOR2X1 _11978_ (
    .A(_05547_),
    .B(_05548_),
    .Y(_05550_)
  );
  NAND2X1 _11979_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05118_),
    .Y(_05551_)
  );
  NOR2X1 _11980_ (
    .A(_05059_),
    .B(_05125_),
    .Y(_05552_)
  );
  NOR2X1 _11981_ (
    .A(_05059_),
    .B(_05121_),
    .Y(_05553_)
  );
  NAND2X1 _11982_ (
    .A(_05508_),
    .B(_05552_),
    .Y(_05554_)
  );
  XNOR2X1 _11983_ (
    .A(_05508_),
    .B(_05552_),
    .Y(_05555_)
  );
  XOR2X1 _11984_ (
    .A(_05551_),
    .B(_05555_),
    .Y(_05556_)
  );
  AOI21X1 _11985_ (
    .A(_05550_),
    .B(_05556_),
    .C(_05549_),
    .Y(_05557_)
  );
  XNOR2X1 _11986_ (
    .A(_05505_),
    .B(_05511_),
    .Y(_05558_)
  );
  NOR2X1 _11987_ (
    .A(_05557_),
    .B(_05558_),
    .Y(_05559_)
  );
  XOR2X1 _11988_ (
    .A(_05557_),
    .B(_05558_),
    .Y(_05560_)
  );
  NAND2X1 _11989_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05164_),
    .Y(_05561_)
  );
  AND2X1 _11990_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05159_),
    .Y(_05562_)
  );
  NAND3X1 _11991_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05164_),
    .C(_05517_),
    .Y(_05563_)
  );
  XOR2X1 _11992_ (
    .A(_05517_),
    .B(_05561_),
    .Y(_05564_)
  );
  NAND2X1 _11993_ (
    .A(multiplier_0.op1_11_ ),
    .B(_05169_),
    .Y(_05565_)
  );
  OAI21X1 _11994_ (
    .A(_05564_),
    .B(_05565_),
    .C(_05563_),
    .Y(_05566_)
  );
  XOR2X1 _11995_ (
    .A(_05519_),
    .B(_05520_),
    .Y(_05567_)
  );
  OAI21X1 _11996_ (
    .A(_05551_),
    .B(_05555_),
    .C(_05554_),
    .Y(_05568_)
  );
  NAND2X1 _11997_ (
    .A(_05567_),
    .B(_05568_),
    .Y(_05569_)
  );
  XOR2X1 _11998_ (
    .A(_05567_),
    .B(_05568_),
    .Y(_05570_)
  );
  NAND2X1 _11999_ (
    .A(_05566_),
    .B(_05570_),
    .Y(_05571_)
  );
  XOR2X1 _12000_ (
    .A(_05566_),
    .B(_05570_),
    .Y(_05572_)
  );
  AOI21X1 _12001_ (
    .A(_05560_),
    .B(_05572_),
    .C(_05559_),
    .Y(_05573_)
  );
  XNOR2X1 _12002_ (
    .A(_05515_),
    .B(_05527_),
    .Y(_05574_)
  );
  OR2X1 _12003_ (
    .A(_05573_),
    .B(_05574_),
    .Y(_05575_)
  );
  NAND2X1 _12004_ (
    .A(_05569_),
    .B(_05571_),
    .Y(_05576_)
  );
  XOR2X1 _12005_ (
    .A(_05573_),
    .B(_05574_),
    .Y(_05577_)
  );
  NAND2X1 _12006_ (
    .A(_05576_),
    .B(_05577_),
    .Y(_05578_)
  );
  OAI21X1 _12007_ (
    .A(_05573_),
    .B(_05574_),
    .C(_05578_),
    .Y(_05579_)
  );
  XNOR2X1 _12008_ (
    .A(_05531_),
    .B(_05532_),
    .Y(_05580_)
  );
  AOI21X1 _12009_ (
    .A(_05575_),
    .B(_05578_),
    .C(_05580_),
    .Y(_05581_)
  );
  XNOR2X1 _12010_ (
    .A(_05534_),
    .B(_05535_),
    .Y(_05582_)
  );
  NAND2X1 _12011_ (
    .A(_05581_),
    .B(_05582_),
    .Y(_05583_)
  );
  AND2X1 _12012_ (
    .A(multiplier_0.op1_2_ ),
    .B(_05098_),
    .Y(_05584_)
  );
  NOR2X1 _12013_ (
    .A(multiplier_0.op1_1_ ),
    .B(_05100_),
    .Y(_05585_)
  );
  NAND2X1 _12014_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05104_),
    .Y(_05586_)
  );
  XNOR2X1 _12015_ (
    .A(_05584_),
    .B(_05585_),
    .Y(_05587_)
  );
  NOR2X1 _12016_ (
    .A(_05586_),
    .B(_05587_),
    .Y(_05588_)
  );
  AOI21X1 _12017_ (
    .A(_05584_),
    .B(_05585_),
    .C(_05588_),
    .Y(_05589_)
  );
  XNOR2X1 _12018_ (
    .A(_05544_),
    .B(_05545_),
    .Y(_05590_)
  );
  NOR2X1 _12019_ (
    .A(_05589_),
    .B(_05590_),
    .Y(_05591_)
  );
  XOR2X1 _12020_ (
    .A(_05589_),
    .B(_05590_),
    .Y(_05592_)
  );
  NAND2X1 _12021_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05118_),
    .Y(_05593_)
  );
  NAND2X1 _12022_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05126_),
    .Y(_05594_)
  );
  NAND3X1 _12023_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05126_),
    .C(_05553_),
    .Y(_05595_)
  );
  XOR2X1 _12024_ (
    .A(_05553_),
    .B(_05594_),
    .Y(_05596_)
  );
  XOR2X1 _12025_ (
    .A(_05593_),
    .B(_05596_),
    .Y(_05597_)
  );
  AOI21X1 _12026_ (
    .A(_05592_),
    .B(_05597_),
    .C(_05591_),
    .Y(_05598_)
  );
  XNOR2X1 _12027_ (
    .A(_05550_),
    .B(_05556_),
    .Y(_05599_)
  );
  NOR2X1 _12028_ (
    .A(_05598_),
    .B(_05599_),
    .Y(_05600_)
  );
  XOR2X1 _12029_ (
    .A(_05598_),
    .B(_05599_),
    .Y(_05601_)
  );
  NAND2X1 _12030_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05164_),
    .Y(_05602_)
  );
  NAND3X1 _12031_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05164_),
    .C(_05562_),
    .Y(_05603_)
  );
  XOR2X1 _12032_ (
    .A(_05562_),
    .B(_05602_),
    .Y(_05604_)
  );
  NAND2X1 _12033_ (
    .A(multiplier_0.op1_10_ ),
    .B(_05169_),
    .Y(_05605_)
  );
  OAI21X1 _12034_ (
    .A(_05604_),
    .B(_05605_),
    .C(_05603_),
    .Y(_05606_)
  );
  XOR2X1 _12035_ (
    .A(_05564_),
    .B(_05565_),
    .Y(_05607_)
  );
  OAI21X1 _12036_ (
    .A(_05593_),
    .B(_05596_),
    .C(_05595_),
    .Y(_05608_)
  );
  NAND2X1 _12037_ (
    .A(_05607_),
    .B(_05608_),
    .Y(_05609_)
  );
  XOR2X1 _12038_ (
    .A(_05607_),
    .B(_05608_),
    .Y(_05610_)
  );
  NAND2X1 _12039_ (
    .A(_05606_),
    .B(_05610_),
    .Y(_05611_)
  );
  XNOR2X1 _12040_ (
    .A(_05606_),
    .B(_05610_),
    .Y(_05612_)
  );
  INVX1 _12041_ (
    .A(_05612_),
    .Y(_05613_)
  );
  AOI21X1 _12042_ (
    .A(_05601_),
    .B(_05613_),
    .C(_05600_),
    .Y(_05614_)
  );
  XNOR2X1 _12043_ (
    .A(_05560_),
    .B(_05572_),
    .Y(_05615_)
  );
  OR2X1 _12044_ (
    .A(_05614_),
    .B(_05615_),
    .Y(_05616_)
  );
  NAND2X1 _12045_ (
    .A(_05609_),
    .B(_05611_),
    .Y(_05617_)
  );
  XOR2X1 _12046_ (
    .A(_05614_),
    .B(_05615_),
    .Y(_05618_)
  );
  NAND2X1 _12047_ (
    .A(_05617_),
    .B(_05618_),
    .Y(_05619_)
  );
  OAI21X1 _12048_ (
    .A(_05614_),
    .B(_05615_),
    .C(_05619_),
    .Y(_05620_)
  );
  XNOR2X1 _12049_ (
    .A(_05576_),
    .B(_05577_),
    .Y(_05621_)
  );
  AOI21X1 _12050_ (
    .A(_05616_),
    .B(_05619_),
    .C(_05621_),
    .Y(_05622_)
  );
  XNOR2X1 _12051_ (
    .A(_05579_),
    .B(_05580_),
    .Y(_05623_)
  );
  AND2X1 _12052_ (
    .A(_05622_),
    .B(_05623_),
    .Y(_05624_)
  );
  XNOR2X1 _12053_ (
    .A(_05622_),
    .B(_05623_),
    .Y(_05625_)
  );
  INVX1 _12054_ (
    .A(_05625_),
    .Y(_05626_)
  );
  NAND2X1 _12055_ (
    .A(multiplier_0.op1_1_ ),
    .B(_05098_),
    .Y(_05627_)
  );
  AOI21X1 _12056_ (
    .A(multiplier_0.op1_1_ ),
    .B(_05098_),
    .C(_05065_),
    .Y(_05628_)
  );
  OR2X1 _12057_ (
    .A(_05100_),
    .B(_05628_),
    .Y(_05629_)
  );
  XNOR2X1 _12058_ (
    .A(_05586_),
    .B(_05587_),
    .Y(_05630_)
  );
  NOR2X1 _12059_ (
    .A(_05629_),
    .B(_05630_),
    .Y(_05631_)
  );
  XOR2X1 _12060_ (
    .A(_05629_),
    .B(_05630_),
    .Y(_05632_)
  );
  NAND2X1 _12061_ (
    .A(multiplier_0.op1_6_ ),
    .B(_05118_),
    .Y(_05633_)
  );
  NAND2X1 _12062_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05122_),
    .Y(_05634_)
  );
  OAI22X1 _12063_ (
    .A(_05060_),
    .B(_05121_),
    .C(_05125_),
    .D(_05061_),
    .Y(_05635_)
  );
  OAI21X1 _12064_ (
    .A(_05594_),
    .B(_05634_),
    .C(_05635_),
    .Y(_05636_)
  );
  XNOR2X1 _12065_ (
    .A(_05633_),
    .B(_05636_),
    .Y(_05637_)
  );
  INVX1 _12066_ (
    .A(_05637_),
    .Y(_05638_)
  );
  AOI21X1 _12067_ (
    .A(_05632_),
    .B(_05638_),
    .C(_05631_),
    .Y(_05639_)
  );
  XNOR2X1 _12068_ (
    .A(_05592_),
    .B(_05597_),
    .Y(_05640_)
  );
  NOR2X1 _12069_ (
    .A(_05639_),
    .B(_05640_),
    .Y(_05641_)
  );
  XOR2X1 _12070_ (
    .A(_05639_),
    .B(_05640_),
    .Y(_05642_)
  );
  NAND2X1 _12071_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05159_),
    .Y(_05643_)
  );
  NOR2X1 _12072_ (
    .A(_05602_),
    .B(_05643_),
    .Y(_05644_)
  );
  AOI22X1 _12073_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05159_),
    .C(_05164_),
    .D(multiplier_0.op1_7_ ),
    .Y(_05645_)
  );
  OR2X1 _12074_ (
    .A(_05644_),
    .B(_05645_),
    .Y(_05646_)
  );
  NAND2X1 _12075_ (
    .A(multiplier_0.op1_9_ ),
    .B(_05169_),
    .Y(_05647_)
  );
  NOR2X1 _12076_ (
    .A(_05646_),
    .B(_05647_),
    .Y(_05648_)
  );
  NOR2X1 _12077_ (
    .A(_05644_),
    .B(_05648_),
    .Y(_05649_)
  );
  XOR2X1 _12078_ (
    .A(_05604_),
    .B(_05605_),
    .Y(_05650_)
  );
  OAI22X1 _12079_ (
    .A(_05594_),
    .B(_05634_),
    .C(_05636_),
    .D(_05633_),
    .Y(_05651_)
  );
  NAND2X1 _12080_ (
    .A(_05650_),
    .B(_05651_),
    .Y(_05652_)
  );
  XOR2X1 _12081_ (
    .A(_05650_),
    .B(_05651_),
    .Y(_05653_)
  );
  OAI21X1 _12082_ (
    .A(_05644_),
    .B(_05648_),
    .C(_05653_),
    .Y(_05654_)
  );
  XNOR2X1 _12083_ (
    .A(_05649_),
    .B(_05653_),
    .Y(_05655_)
  );
  AOI21X1 _12084_ (
    .A(_05642_),
    .B(_05655_),
    .C(_05641_),
    .Y(_05656_)
  );
  XNOR2X1 _12085_ (
    .A(_05601_),
    .B(_05613_),
    .Y(_05657_)
  );
  OR2X1 _12086_ (
    .A(_05656_),
    .B(_05657_),
    .Y(_05658_)
  );
  NAND2X1 _12087_ (
    .A(_05652_),
    .B(_05654_),
    .Y(_05659_)
  );
  XOR2X1 _12088_ (
    .A(_05656_),
    .B(_05657_),
    .Y(_05660_)
  );
  NAND2X1 _12089_ (
    .A(_05659_),
    .B(_05660_),
    .Y(_05661_)
  );
  OAI21X1 _12090_ (
    .A(_05656_),
    .B(_05657_),
    .C(_05661_),
    .Y(_05662_)
  );
  XNOR2X1 _12091_ (
    .A(_05617_),
    .B(_05618_),
    .Y(_05663_)
  );
  AOI21X1 _12092_ (
    .A(_05658_),
    .B(_05661_),
    .C(_05663_),
    .Y(_05664_)
  );
  XNOR2X1 _12093_ (
    .A(_05620_),
    .B(_05621_),
    .Y(_05665_)
  );
  NAND2X1 _12094_ (
    .A(_05664_),
    .B(_05665_),
    .Y(_05666_)
  );
  XNOR2X1 _12095_ (
    .A(_05664_),
    .B(_05665_),
    .Y(_05667_)
  );
  NAND2X1 _12096_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05098_),
    .Y(_05668_)
  );
  NAND2X1 _12097_ (
    .A(multiplier_0.op1_1_ ),
    .B(_05104_),
    .Y(_05669_)
  );
  NAND2X1 _12098_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05104_),
    .Y(_05670_)
  );
  NOR2X1 _12099_ (
    .A(_05627_),
    .B(_05670_),
    .Y(_05671_)
  );
  OAI21X1 _12100_ (
    .A(_05049_),
    .B(_05097_),
    .C(_05671_),
    .Y(_05672_)
  );
  NAND2X1 _12101_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05126_),
    .Y(_05673_)
  );
  NAND2X1 _12102_ (
    .A(multiplier_0.op1_2_ ),
    .B(_05104_),
    .Y(_05674_)
  );
  NOR2X1 _12103_ (
    .A(_05063_),
    .B(_05125_),
    .Y(_05675_)
  );
  OR2X1 _12104_ (
    .A(_05673_),
    .B(_05674_),
    .Y(_05676_)
  );
  XNOR2X1 _12105_ (
    .A(_05673_),
    .B(_05674_),
    .Y(_05677_)
  );
  XNOR2X1 _12106_ (
    .A(_05634_),
    .B(_05677_),
    .Y(_05678_)
  );
  NOR2X1 _12107_ (
    .A(_05065_),
    .B(_05100_),
    .Y(_05679_)
  );
  AOI21X1 _12108_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05104_),
    .C(_05627_),
    .Y(_05680_)
  );
  XNOR2X1 _12109_ (
    .A(_05679_),
    .B(_05680_),
    .Y(_05681_)
  );
  OAI21X1 _12110_ (
    .A(_05678_),
    .B(_05681_),
    .C(_05672_),
    .Y(_05682_)
  );
  XNOR2X1 _12111_ (
    .A(_05632_),
    .B(_05638_),
    .Y(_05683_)
  );
  INVX1 _12112_ (
    .A(_05683_),
    .Y(_05684_)
  );
  NAND2X1 _12113_ (
    .A(_05682_),
    .B(_05684_),
    .Y(_05685_)
  );
  XOR2X1 _12114_ (
    .A(_05682_),
    .B(_05683_),
    .Y(_05686_)
  );
  NAND2X1 _12115_ (
    .A(multiplier_0.op1_6_ ),
    .B(_05164_),
    .Y(_05687_)
  );
  NAND2X1 _12116_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05118_),
    .Y(_05688_)
  );
  NOR2X1 _12117_ (
    .A(_05060_),
    .B(_05163_),
    .Y(_05689_)
  );
  OR2X1 _12118_ (
    .A(_05060_),
    .B(_05163_),
    .Y(_05690_)
  );
  XNOR2X1 _12119_ (
    .A(_05687_),
    .B(_05688_),
    .Y(_05691_)
  );
  OAI22X1 _12120_ (
    .A(_05633_),
    .B(_05690_),
    .C(_05691_),
    .D(_05643_),
    .Y(_05692_)
  );
  XOR2X1 _12121_ (
    .A(_05646_),
    .B(_05647_),
    .Y(_05693_)
  );
  OAI21X1 _12122_ (
    .A(_05634_),
    .B(_05677_),
    .C(_05676_),
    .Y(_05694_)
  );
  NAND2X1 _12123_ (
    .A(_05693_),
    .B(_05694_),
    .Y(_05695_)
  );
  XOR2X1 _12124_ (
    .A(_05693_),
    .B(_05694_),
    .Y(_05696_)
  );
  NAND2X1 _12125_ (
    .A(_05692_),
    .B(_05696_),
    .Y(_05697_)
  );
  XNOR2X1 _12126_ (
    .A(_05692_),
    .B(_05696_),
    .Y(_05698_)
  );
  OAI21X1 _12127_ (
    .A(_05686_),
    .B(_05698_),
    .C(_05685_),
    .Y(_05699_)
  );
  XNOR2X1 _12128_ (
    .A(_05642_),
    .B(_05655_),
    .Y(_05700_)
  );
  INVX1 _12129_ (
    .A(_05700_),
    .Y(_05701_)
  );
  NAND2X1 _12130_ (
    .A(_05699_),
    .B(_05701_),
    .Y(_05702_)
  );
  NAND2X1 _12131_ (
    .A(_05695_),
    .B(_05697_),
    .Y(_05703_)
  );
  XOR2X1 _12132_ (
    .A(_05699_),
    .B(_05700_),
    .Y(_05704_)
  );
  INVX1 _12133_ (
    .A(_05704_),
    .Y(_05705_)
  );
  NAND2X1 _12134_ (
    .A(_05703_),
    .B(_05705_),
    .Y(_05706_)
  );
  NAND2X1 _12135_ (
    .A(_05702_),
    .B(_05706_),
    .Y(_05707_)
  );
  XNOR2X1 _12136_ (
    .A(_05659_),
    .B(_05660_),
    .Y(_05708_)
  );
  AOI21X1 _12137_ (
    .A(_05702_),
    .B(_05706_),
    .C(_05708_),
    .Y(_05709_)
  );
  XNOR2X1 _12138_ (
    .A(_05662_),
    .B(_05663_),
    .Y(_05710_)
  );
  AND2X1 _12139_ (
    .A(_05709_),
    .B(_05710_),
    .Y(_05711_)
  );
  NOR2X1 _12140_ (
    .A(_05709_),
    .B(_05710_),
    .Y(_05712_)
  );
  NOR2X1 _12141_ (
    .A(_05711_),
    .B(_05712_),
    .Y(_05713_)
  );
  XNOR2X1 _12142_ (
    .A(_05668_),
    .B(_05669_),
    .Y(_05714_)
  );
  NAND2X1 _12143_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05118_),
    .Y(_05715_)
  );
  NOR2X1 _12144_ (
    .A(_05062_),
    .B(_05121_),
    .Y(_05716_)
  );
  NOR2X1 _12145_ (
    .A(_05063_),
    .B(_05121_),
    .Y(_05717_)
  );
  NAND2X1 _12146_ (
    .A(_05675_),
    .B(_05716_),
    .Y(_05718_)
  );
  XNOR2X1 _12147_ (
    .A(_05675_),
    .B(_05716_),
    .Y(_05719_)
  );
  XNOR2X1 _12148_ (
    .A(_05715_),
    .B(_05719_),
    .Y(_05720_)
  );
  NOR2X1 _12149_ (
    .A(_05714_),
    .B(_05720_),
    .Y(_05721_)
  );
  XNOR2X1 _12150_ (
    .A(_05678_),
    .B(_05681_),
    .Y(_05722_)
  );
  INVX1 _12151_ (
    .A(_05722_),
    .Y(_05723_)
  );
  NAND2X1 _12152_ (
    .A(_05721_),
    .B(_05723_),
    .Y(_05724_)
  );
  XOR2X1 _12153_ (
    .A(_05721_),
    .B(_05722_),
    .Y(_05725_)
  );
  NOR2X1 _12154_ (
    .A(_05059_),
    .B(_05158_),
    .Y(_05726_)
  );
  NAND2X1 _12155_ (
    .A(_05689_),
    .B(_05726_),
    .Y(_05727_)
  );
  NOR2X1 _12156_ (
    .A(_05689_),
    .B(_05726_),
    .Y(_05728_)
  );
  XNOR2X1 _12157_ (
    .A(_05690_),
    .B(_05726_),
    .Y(_05729_)
  );
  NAND2X1 _12158_ (
    .A(multiplier_0.op1_7_ ),
    .B(_05169_),
    .Y(_05730_)
  );
  OAI21X1 _12159_ (
    .A(_05728_),
    .B(_05730_),
    .C(_05727_),
    .Y(_05731_)
  );
  XNOR2X1 _12160_ (
    .A(_05643_),
    .B(_05691_),
    .Y(_05732_)
  );
  OAI21X1 _12161_ (
    .A(_05715_),
    .B(_05719_),
    .C(_05718_),
    .Y(_05733_)
  );
  INVX1 _12162_ (
    .A(_05733_),
    .Y(_05734_)
  );
  XNOR2X1 _12163_ (
    .A(_05732_),
    .B(_05734_),
    .Y(_05735_)
  );
  INVX1 _12164_ (
    .A(_05735_),
    .Y(_05736_)
  );
  NAND2X1 _12165_ (
    .A(_05731_),
    .B(_05736_),
    .Y(_05737_)
  );
  XOR2X1 _12166_ (
    .A(_05731_),
    .B(_05735_),
    .Y(_05738_)
  );
  OAI21X1 _12167_ (
    .A(_05725_),
    .B(_05738_),
    .C(_05724_),
    .Y(_05739_)
  );
  XOR2X1 _12168_ (
    .A(_05686_),
    .B(_05698_),
    .Y(_05740_)
  );
  NAND2X1 _12169_ (
    .A(_05739_),
    .B(_05740_),
    .Y(_05741_)
  );
  OAI21X1 _12170_ (
    .A(_05732_),
    .B(_05734_),
    .C(_05737_),
    .Y(_05742_)
  );
  INVX1 _12171_ (
    .A(_05742_),
    .Y(_05743_)
  );
  XNOR2X1 _12172_ (
    .A(_05739_),
    .B(_05740_),
    .Y(_05744_)
  );
  OAI21X1 _12173_ (
    .A(_05743_),
    .B(_05744_),
    .C(_05741_),
    .Y(_05745_)
  );
  XNOR2X1 _12174_ (
    .A(_05703_),
    .B(_05704_),
    .Y(_05746_)
  );
  NAND2X1 _12175_ (
    .A(_05745_),
    .B(_05746_),
    .Y(_05747_)
  );
  XOR2X1 _12176_ (
    .A(_05707_),
    .B(_05708_),
    .Y(_05748_)
  );
  OR2X1 _12177_ (
    .A(_05747_),
    .B(_05748_),
    .Y(_05749_)
  );
  XNOR2X1 _12178_ (
    .A(_05747_),
    .B(_05748_),
    .Y(_05750_)
  );
  NAND2X1 _12179_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05118_),
    .Y(_05751_)
  );
  NOR2X1 _12180_ (
    .A(_05064_),
    .B(_05125_),
    .Y(_05752_)
  );
  NOR2X1 _12181_ (
    .A(_05064_),
    .B(_05121_),
    .Y(_05753_)
  );
  NAND2X1 _12182_ (
    .A(multiplier_0.op1_1_ ),
    .B(_05122_),
    .Y(_05754_)
  );
  NAND2X1 _12183_ (
    .A(_05675_),
    .B(_05753_),
    .Y(_05755_)
  );
  XNOR2X1 _12184_ (
    .A(_05717_),
    .B(_05752_),
    .Y(_05756_)
  );
  XNOR2X1 _12185_ (
    .A(_05751_),
    .B(_05756_),
    .Y(_05757_)
  );
  NOR2X1 _12186_ (
    .A(_05670_),
    .B(_05757_),
    .Y(_05758_)
  );
  XOR2X1 _12187_ (
    .A(_05714_),
    .B(_05720_),
    .Y(_05759_)
  );
  NAND2X1 _12188_ (
    .A(_05758_),
    .B(_05759_),
    .Y(_05760_)
  );
  XNOR2X1 _12189_ (
    .A(_05758_),
    .B(_05759_),
    .Y(_05761_)
  );
  NOR2X1 _12190_ (
    .A(_05061_),
    .B(_05163_),
    .Y(_05762_)
  );
  OR2X1 _12191_ (
    .A(_05061_),
    .B(_05158_),
    .Y(_05763_)
  );
  OAI22X1 _12192_ (
    .A(_05060_),
    .B(_05158_),
    .C(_05163_),
    .D(_05061_),
    .Y(_05764_)
  );
  OAI21X1 _12193_ (
    .A(_05690_),
    .B(_05763_),
    .C(_05764_),
    .Y(_05765_)
  );
  NAND2X1 _12194_ (
    .A(multiplier_0.op1_6_ ),
    .B(_05169_),
    .Y(_05766_)
  );
  OAI22X1 _12195_ (
    .A(_05690_),
    .B(_05763_),
    .C(_05765_),
    .D(_05766_),
    .Y(_05767_)
  );
  XNOR2X1 _12196_ (
    .A(_05729_),
    .B(_05730_),
    .Y(_05768_)
  );
  OAI21X1 _12197_ (
    .A(_05751_),
    .B(_05756_),
    .C(_05755_),
    .Y(_05769_)
  );
  NAND2X1 _12198_ (
    .A(_05768_),
    .B(_05769_),
    .Y(_05770_)
  );
  XOR2X1 _12199_ (
    .A(_05768_),
    .B(_05769_),
    .Y(_05771_)
  );
  NAND2X1 _12200_ (
    .A(_05767_),
    .B(_05771_),
    .Y(_05772_)
  );
  XNOR2X1 _12201_ (
    .A(_05767_),
    .B(_05771_),
    .Y(_05773_)
  );
  OAI21X1 _12202_ (
    .A(_05761_),
    .B(_05773_),
    .C(_05760_),
    .Y(_05774_)
  );
  XOR2X1 _12203_ (
    .A(_05725_),
    .B(_05738_),
    .Y(_05775_)
  );
  NAND2X1 _12204_ (
    .A(_05774_),
    .B(_05775_),
    .Y(_05776_)
  );
  XNOR2X1 _12205_ (
    .A(_05774_),
    .B(_05775_),
    .Y(_05777_)
  );
  INVX1 _12206_ (
    .A(_05777_),
    .Y(_05778_)
  );
  NAND2X1 _12207_ (
    .A(_05770_),
    .B(_05772_),
    .Y(_05779_)
  );
  NAND2X1 _12208_ (
    .A(_05778_),
    .B(_05779_),
    .Y(_05780_)
  );
  NAND2X1 _12209_ (
    .A(_05776_),
    .B(_05780_),
    .Y(_05781_)
  );
  XNOR2X1 _12210_ (
    .A(_05743_),
    .B(_05744_),
    .Y(_05782_)
  );
  INVX1 _12211_ (
    .A(_05782_),
    .Y(_05783_)
  );
  NAND2X1 _12212_ (
    .A(_05781_),
    .B(_05783_),
    .Y(_05784_)
  );
  XNOR2X1 _12213_ (
    .A(_05745_),
    .B(_05746_),
    .Y(_05785_)
  );
  NOR2X1 _12214_ (
    .A(_05784_),
    .B(_05785_),
    .Y(_05786_)
  );
  XOR2X1 _12215_ (
    .A(_05784_),
    .B(_05785_),
    .Y(_05787_)
  );
  XNOR2X1 _12216_ (
    .A(_05670_),
    .B(_05757_),
    .Y(_05788_)
  );
  NOR2X1 _12217_ (
    .A(_05062_),
    .B(_05163_),
    .Y(_05789_)
  );
  NOR2X1 _12218_ (
    .A(_05062_),
    .B(_05158_),
    .Y(_05790_)
  );
  XOR2X1 _12219_ (
    .A(_05763_),
    .B(_05789_),
    .Y(_05791_)
  );
  NAND2X1 _12220_ (
    .A(multiplier_0.op1_5_ ),
    .B(_05169_),
    .Y(_05792_)
  );
  NOR2X1 _12221_ (
    .A(_05791_),
    .B(_05792_),
    .Y(_05793_)
  );
  AOI21X1 _12222_ (
    .A(_05762_),
    .B(_05790_),
    .C(_05793_),
    .Y(_05794_)
  );
  XOR2X1 _12223_ (
    .A(_05765_),
    .B(_05766_),
    .Y(_05795_)
  );
  NOR2X1 _12224_ (
    .A(_05065_),
    .B(_05121_),
    .Y(_05796_)
  );
  NAND2X1 _12225_ (
    .A(_05752_),
    .B(_05796_),
    .Y(_05797_)
  );
  AOI21X1 _12226_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05126_),
    .C(_05753_),
    .Y(_05798_)
  );
  AOI21X1 _12227_ (
    .A(_05752_),
    .B(_05796_),
    .C(_05798_),
    .Y(_05799_)
  );
  NAND2X1 _12228_ (
    .A(multiplier_0.op1_2_ ),
    .B(_05118_),
    .Y(_05800_)
  );
  OAI21X1 _12229_ (
    .A(_05798_),
    .B(_05800_),
    .C(_05797_),
    .Y(_05801_)
  );
  NAND2X1 _12230_ (
    .A(_05795_),
    .B(_05801_),
    .Y(_05802_)
  );
  NOR2X1 _12231_ (
    .A(_05795_),
    .B(_05801_),
    .Y(_05803_)
  );
  XNOR2X1 _12232_ (
    .A(_05795_),
    .B(_05801_),
    .Y(_05804_)
  );
  XNOR2X1 _12233_ (
    .A(_05794_),
    .B(_05804_),
    .Y(_05805_)
  );
  NOR2X1 _12234_ (
    .A(_05788_),
    .B(_05805_),
    .Y(_05806_)
  );
  XOR2X1 _12235_ (
    .A(_05761_),
    .B(_05773_),
    .Y(_05807_)
  );
  NAND2X1 _12236_ (
    .A(_05806_),
    .B(_05807_),
    .Y(_05808_)
  );
  OAI21X1 _12237_ (
    .A(_05794_),
    .B(_05803_),
    .C(_05802_),
    .Y(_05809_)
  );
  INVX1 _12238_ (
    .A(_05809_),
    .Y(_05810_)
  );
  XNOR2X1 _12239_ (
    .A(_05806_),
    .B(_05807_),
    .Y(_05811_)
  );
  OAI21X1 _12240_ (
    .A(_05810_),
    .B(_05811_),
    .C(_05808_),
    .Y(_05812_)
  );
  INVX1 _12241_ (
    .A(_05812_),
    .Y(_05813_)
  );
  XOR2X1 _12242_ (
    .A(_05777_),
    .B(_05779_),
    .Y(_05814_)
  );
  NOR2X1 _12243_ (
    .A(_05813_),
    .B(_05814_),
    .Y(_05815_)
  );
  NAND2X1 _12244_ (
    .A(multiplier_0.op1_8_ ),
    .B(_05169_),
    .Y(_05816_)
  );
  XNOR2X1 _12245_ (
    .A(_05813_),
    .B(_05814_),
    .Y(_05817_)
  );
  NOR2X1 _12246_ (
    .A(_05816_),
    .B(_05817_),
    .Y(_05818_)
  );
  NOR2X1 _12247_ (
    .A(_05815_),
    .B(_05818_),
    .Y(_05819_)
  );
  XNOR2X1 _12248_ (
    .A(_05781_),
    .B(_05783_),
    .Y(_05820_)
  );
  OR2X1 _12249_ (
    .A(_05819_),
    .B(_05820_),
    .Y(_05821_)
  );
  XNOR2X1 _12250_ (
    .A(_05799_),
    .B(_05800_),
    .Y(_05822_)
  );
  INVX1 _12251_ (
    .A(_05822_),
    .Y(_05823_)
  );
  OR2X1 _12252_ (
    .A(_05063_),
    .B(_05163_),
    .Y(_05824_)
  );
  NAND3X1 _12253_ (
    .A(multiplier_0.op1_2_ ),
    .B(_05164_),
    .C(_05790_),
    .Y(_05825_)
  );
  XOR2X1 _12254_ (
    .A(_05790_),
    .B(_05824_),
    .Y(_05826_)
  );
  NAND2X1 _12255_ (
    .A(multiplier_0.op1_4_ ),
    .B(_05169_),
    .Y(_05827_)
  );
  OAI21X1 _12256_ (
    .A(_05826_),
    .B(_05827_),
    .C(_05825_),
    .Y(_05828_)
  );
  NAND2X1 _12257_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05118_),
    .Y(_05829_)
  );
  NOR2X1 _12258_ (
    .A(_05754_),
    .B(_05829_),
    .Y(_05830_)
  );
  XOR2X1 _12259_ (
    .A(_05791_),
    .B(_05792_),
    .Y(_05831_)
  );
  NAND2X1 _12260_ (
    .A(_05830_),
    .B(_05831_),
    .Y(_05832_)
  );
  XOR2X1 _12261_ (
    .A(_05830_),
    .B(_05831_),
    .Y(_05833_)
  );
  NAND2X1 _12262_ (
    .A(_05828_),
    .B(_05833_),
    .Y(_05834_)
  );
  XNOR2X1 _12263_ (
    .A(_05828_),
    .B(_05833_),
    .Y(_05835_)
  );
  NOR2X1 _12264_ (
    .A(_05823_),
    .B(_05835_),
    .Y(_05836_)
  );
  XOR2X1 _12265_ (
    .A(_05788_),
    .B(_05805_),
    .Y(_05837_)
  );
  AND2X1 _12266_ (
    .A(_05836_),
    .B(_05837_),
    .Y(_05838_)
  );
  XNOR2X1 _12267_ (
    .A(_05836_),
    .B(_05837_),
    .Y(_05839_)
  );
  NAND2X1 _12268_ (
    .A(_05832_),
    .B(_05834_),
    .Y(_05840_)
  );
  AOI21X1 _12269_ (
    .A(_05832_),
    .B(_05834_),
    .C(_05839_),
    .Y(_05841_)
  );
  NOR2X1 _12270_ (
    .A(_05838_),
    .B(_05841_),
    .Y(_05842_)
  );
  XNOR2X1 _12271_ (
    .A(_05809_),
    .B(_05811_),
    .Y(_05843_)
  );
  OAI21X1 _12272_ (
    .A(_05838_),
    .B(_05841_),
    .C(_05843_),
    .Y(_05844_)
  );
  XNOR2X1 _12273_ (
    .A(_05816_),
    .B(_05817_),
    .Y(_05845_)
  );
  NOR2X1 _12274_ (
    .A(_05844_),
    .B(_05845_),
    .Y(_05846_)
  );
  XOR2X1 _12275_ (
    .A(_05839_),
    .B(_05840_),
    .Y(_05847_)
  );
  XNOR2X1 _12276_ (
    .A(_05822_),
    .B(_05835_),
    .Y(_05848_)
  );
  NOR2X1 _12277_ (
    .A(_05064_),
    .B(_05158_),
    .Y(_04442_)
  );
  OR2X1 _12278_ (
    .A(_05064_),
    .B(_05158_),
    .Y(_04443_)
  );
  OAI22X1 _12279_ (
    .A(_05063_),
    .B(_05158_),
    .C(_05163_),
    .D(_05064_),
    .Y(_04444_)
  );
  OAI21X1 _12280_ (
    .A(_05824_),
    .B(_04443_),
    .C(_04444_),
    .Y(_04445_)
  );
  NAND2X1 _12281_ (
    .A(multiplier_0.op1_3_ ),
    .B(_05169_),
    .Y(_04446_)
  );
  OAI22X1 _12282_ (
    .A(_05824_),
    .B(_04443_),
    .C(_04445_),
    .D(_04446_),
    .Y(_04447_)
  );
  XOR2X1 _12283_ (
    .A(_05826_),
    .B(_05827_),
    .Y(_04448_)
  );
  NAND2X1 _12284_ (
    .A(_04447_),
    .B(_04448_),
    .Y(_04449_)
  );
  AOI21X1 _12285_ (
    .A(multiplier_0.op1_1_ ),
    .B(_05118_),
    .C(_05796_),
    .Y(_04450_)
  );
  OR2X1 _12286_ (
    .A(_05830_),
    .B(_04450_),
    .Y(_04451_)
  );
  XNOR2X1 _12287_ (
    .A(_04447_),
    .B(_04448_),
    .Y(_04452_)
  );
  OAI21X1 _12288_ (
    .A(_04451_),
    .B(_04452_),
    .C(_04449_),
    .Y(_04453_)
  );
  NAND2X1 _12289_ (
    .A(_05848_),
    .B(_04453_),
    .Y(_04454_)
  );
  OR2X1 _12290_ (
    .A(_05847_),
    .B(_04454_),
    .Y(_04455_)
  );
  XOR2X1 _12291_ (
    .A(_05842_),
    .B(_05843_),
    .Y(_04456_)
  );
  OR2X1 _12292_ (
    .A(_04455_),
    .B(_04456_),
    .Y(_04457_)
  );
  XOR2X1 _12293_ (
    .A(_04451_),
    .B(_04452_),
    .Y(_04458_)
  );
  NOR2X1 _12294_ (
    .A(_05065_),
    .B(_05163_),
    .Y(_04459_)
  );
  NAND2X1 _12295_ (
    .A(_04442_),
    .B(_04459_),
    .Y(_04460_)
  );
  NAND2X1 _12296_ (
    .A(multiplier_0.op1_2_ ),
    .B(_05169_),
    .Y(_04461_)
  );
  XNOR2X1 _12297_ (
    .A(_04442_),
    .B(_04459_),
    .Y(_04462_)
  );
  OAI21X1 _12298_ (
    .A(_04461_),
    .B(_04462_),
    .C(_04460_),
    .Y(_04463_)
  );
  XOR2X1 _12299_ (
    .A(_04445_),
    .B(_04446_),
    .Y(_04464_)
  );
  NAND2X1 _12300_ (
    .A(_04463_),
    .B(_04464_),
    .Y(_04465_)
  );
  XNOR2X1 _12301_ (
    .A(_04463_),
    .B(_04464_),
    .Y(_04466_)
  );
  OAI21X1 _12302_ (
    .A(_05829_),
    .B(_04466_),
    .C(_04465_),
    .Y(_04467_)
  );
  NAND2X1 _12303_ (
    .A(_04458_),
    .B(_04467_),
    .Y(_04468_)
  );
  XNOR2X1 _12304_ (
    .A(_05848_),
    .B(_04453_),
    .Y(_04469_)
  );
  NOR2X1 _12305_ (
    .A(_04468_),
    .B(_04469_),
    .Y(_04470_)
  );
  XOR2X1 _12306_ (
    .A(_05847_),
    .B(_04454_),
    .Y(_04471_)
  );
  AND2X1 _12307_ (
    .A(_04470_),
    .B(_04471_),
    .Y(_04472_)
  );
  NOR2X1 _12308_ (
    .A(_05065_),
    .B(_05168_),
    .Y(_04473_)
  );
  NAND3X1 _12309_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05169_),
    .C(_04442_),
    .Y(_04474_)
  );
  INVX1 _12310_ (
    .A(_04474_),
    .Y(_04475_)
  );
  XNOR2X1 _12311_ (
    .A(_04461_),
    .B(_04462_),
    .Y(_04476_)
  );
  NOR2X1 _12312_ (
    .A(_04474_),
    .B(_04476_),
    .Y(_04477_)
  );
  INVX1 _12313_ (
    .A(_04477_),
    .Y(_04478_)
  );
  XNOR2X1 _12314_ (
    .A(_05829_),
    .B(_04466_),
    .Y(_04479_)
  );
  OR2X1 _12315_ (
    .A(_04478_),
    .B(_04479_),
    .Y(_04480_)
  );
  INVX1 _12316_ (
    .A(_04480_),
    .Y(_04481_)
  );
  XOR2X1 _12317_ (
    .A(_04458_),
    .B(_04467_),
    .Y(_04482_)
  );
  NAND2X1 _12318_ (
    .A(_04481_),
    .B(_04482_),
    .Y(_04483_)
  );
  INVX1 _12319_ (
    .A(_04483_),
    .Y(_04484_)
  );
  XOR2X1 _12320_ (
    .A(_04468_),
    .B(_04469_),
    .Y(_04485_)
  );
  AND2X1 _12321_ (
    .A(_04484_),
    .B(_04485_),
    .Y(_04486_)
  );
  XOR2X1 _12322_ (
    .A(_04470_),
    .B(_04471_),
    .Y(_04487_)
  );
  AOI21X1 _12323_ (
    .A(_04486_),
    .B(_04487_),
    .C(_04472_),
    .Y(_04488_)
  );
  XNOR2X1 _12324_ (
    .A(_04455_),
    .B(_04456_),
    .Y(_04489_)
  );
  OAI21X1 _12325_ (
    .A(_04488_),
    .B(_04489_),
    .C(_04457_),
    .Y(_04490_)
  );
  XOR2X1 _12326_ (
    .A(_05844_),
    .B(_05845_),
    .Y(_04491_)
  );
  AOI21X1 _12327_ (
    .A(_04490_),
    .B(_04491_),
    .C(_05846_),
    .Y(_04492_)
  );
  XNOR2X1 _12328_ (
    .A(_05819_),
    .B(_05820_),
    .Y(_04493_)
  );
  OAI21X1 _12329_ (
    .A(_04492_),
    .B(_04493_),
    .C(_05821_),
    .Y(_04494_)
  );
  AOI21X1 _12330_ (
    .A(_05787_),
    .B(_04494_),
    .C(_05786_),
    .Y(_04495_)
  );
  OAI21X1 _12331_ (
    .A(_05750_),
    .B(_04495_),
    .C(_05749_),
    .Y(_04496_)
  );
  AOI21X1 _12332_ (
    .A(_05713_),
    .B(_04496_),
    .C(_05711_),
    .Y(_04497_)
  );
  OAI21X1 _12333_ (
    .A(_05667_),
    .B(_04497_),
    .C(_05666_),
    .Y(_04498_)
  );
  AOI21X1 _12334_ (
    .A(_05626_),
    .B(_04498_),
    .C(_05624_),
    .Y(_04499_)
  );
  XNOR2X1 _12335_ (
    .A(_05581_),
    .B(_05582_),
    .Y(_04500_)
  );
  OAI21X1 _12336_ (
    .A(_04499_),
    .B(_04500_),
    .C(_05583_),
    .Y(_04501_)
  );
  AOI21X1 _12337_ (
    .A(_05541_),
    .B(_04501_),
    .C(_05539_),
    .Y(_04502_)
  );
  XNOR2X1 _12338_ (
    .A(_05493_),
    .B(_05495_),
    .Y(_04503_)
  );
  OAI21X1 _12339_ (
    .A(_04502_),
    .B(_04503_),
    .C(_05496_),
    .Y(_04504_)
  );
  AOI21X1 _12340_ (
    .A(_05454_),
    .B(_04504_),
    .C(_05453_),
    .Y(_04505_)
  );
  OAI21X1 _12341_ (
    .A(_05409_),
    .B(_04505_),
    .C(_05407_),
    .Y(_04506_)
  );
  XOR2X1 _12342_ (
    .A(_05359_),
    .B(_05360_),
    .Y(_04507_)
  );
  AOI21X1 _12343_ (
    .A(_04506_),
    .B(_04507_),
    .C(_05361_),
    .Y(_04508_)
  );
  XNOR2X1 _12344_ (
    .A(_05314_),
    .B(_05315_),
    .Y(_04509_)
  );
  INVX1 _12345_ (
    .A(_04509_),
    .Y(_04510_)
  );
  OAI21X1 _12346_ (
    .A(_04508_),
    .B(_04510_),
    .C(_05316_),
    .Y(_04511_)
  );
  XOR2X1 _12347_ (
    .A(_05252_),
    .B(_05278_),
    .Y(_04512_)
  );
  AOI21X1 _12348_ (
    .A(_04511_),
    .B(_04512_),
    .C(_05279_),
    .Y(_04513_)
  );
  AOI21X1 _12349_ (
    .A(_05243_),
    .B(_05269_),
    .C(_05267_),
    .Y(_04514_)
  );
  OAI21X1 _12350_ (
    .A(_05096_),
    .B(_05149_),
    .C(_05100_),
    .Y(_04515_)
  );
  AOI22X1 _12351_ (
    .A(_05104_),
    .B(_05148_),
    .C(_05258_),
    .D(_04515_),
    .Y(_04516_)
  );
  MUX2X1 _12352_ (
    .A(_05264_),
    .B(_05263_),
    .S(_05236_),
    .Y(_04517_)
  );
  XNOR2X1 _12353_ (
    .A(_04516_),
    .B(_04517_),
    .Y(_04518_)
  );
  XNOR2X1 _12354_ (
    .A(_05243_),
    .B(_04518_),
    .Y(_04519_)
  );
  XNOR2X1 _12355_ (
    .A(_04514_),
    .B(_04519_),
    .Y(_04520_)
  );
  MUX2X1 _12356_ (
    .A(_05273_),
    .B(_05271_),
    .S(_05275_),
    .Y(_04521_)
  );
  XNOR2X1 _12357_ (
    .A(_04520_),
    .B(_04521_),
    .Y(_04522_)
  );
  XOR2X1 _12358_ (
    .A(_05277_),
    .B(_04522_),
    .Y(_04523_)
  );
  XNOR2X1 _12359_ (
    .A(_04513_),
    .B(_04523_),
    .Y(_04524_)
  );
  INVX1 _12360_ (
    .A(_04524_),
    .Y(_04525_)
  );
  AOI21X1 _12361_ (
    .A(_05047_),
    .B(_05049_),
    .C(_04525_),
    .Y(_04526_)
  );
  XNOR2X1 _12362_ (
    .A(multiplier_0.reshi_15_ ),
    .B(_04526_),
    .Y(_04527_)
  );
  INVX1 _12363_ (
    .A(_04527_),
    .Y(_04528_)
  );
  XNOR2X1 _12364_ (
    .A(_04511_),
    .B(_04512_),
    .Y(_04529_)
  );
  NAND2X1 _12365_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04529_),
    .Y(_04530_)
  );
  NOR2X1 _12366_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04524_),
    .Y(_04531_)
  );
  OAI21X1 _12367_ (
    .A(_05049_),
    .B(_04525_),
    .C(_05047_),
    .Y(_04532_)
  );
  NAND2X1 _12368_ (
    .A(_04530_),
    .B(_04532_),
    .Y(_04533_)
  );
  NAND3X1 _12369_ (
    .A(multiplier_0.reshi_14_ ),
    .B(_04530_),
    .C(_04532_),
    .Y(_04534_)
  );
  XOR2X1 _12370_ (
    .A(multiplier_0.reshi_14_ ),
    .B(_04533_),
    .Y(_04535_)
  );
  XNOR2X1 _12371_ (
    .A(_04508_),
    .B(_04510_),
    .Y(_04536_)
  );
  NAND2X1 _12372_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04536_),
    .Y(_04537_)
  );
  NAND2X1 _12373_ (
    .A(_04532_),
    .B(_04537_),
    .Y(_04538_)
  );
  OR2X1 _12374_ (
    .A(_05066_),
    .B(_04538_),
    .Y(_04539_)
  );
  INVX1 _12375_ (
    .A(_04539_),
    .Y(_04540_)
  );
  NAND2X1 _12376_ (
    .A(_05066_),
    .B(_04538_),
    .Y(_04541_)
  );
  XNOR2X1 _12377_ (
    .A(_04506_),
    .B(_04507_),
    .Y(_04542_)
  );
  NAND2X1 _12378_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04542_),
    .Y(_04543_)
  );
  AND2X1 _12379_ (
    .A(_04532_),
    .B(_04543_),
    .Y(_04544_)
  );
  NAND2X1 _12380_ (
    .A(multiplier_0.reshi_12_ ),
    .B(_04544_),
    .Y(_04545_)
  );
  XNOR2X1 _12381_ (
    .A(multiplier_0.reshi_12_ ),
    .B(_04544_),
    .Y(_04546_)
  );
  XNOR2X1 _12382_ (
    .A(_05409_),
    .B(_04505_),
    .Y(_04547_)
  );
  NAND2X1 _12383_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04547_),
    .Y(_04548_)
  );
  NAND2X1 _12384_ (
    .A(_04532_),
    .B(_04548_),
    .Y(_04549_)
  );
  NAND2X1 _12385_ (
    .A(_05067_),
    .B(_04549_),
    .Y(_04550_)
  );
  OR2X1 _12386_ (
    .A(_05067_),
    .B(_04549_),
    .Y(_04551_)
  );
  INVX1 _12387_ (
    .A(_04551_),
    .Y(_04552_)
  );
  XNOR2X1 _12388_ (
    .A(_05454_),
    .B(_04504_),
    .Y(_04553_)
  );
  NAND2X1 _12389_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04553_),
    .Y(_04554_)
  );
  NAND2X1 _12390_ (
    .A(_04532_),
    .B(_04554_),
    .Y(_04555_)
  );
  NAND3X1 _12391_ (
    .A(multiplier_0.reshi_10_ ),
    .B(_04532_),
    .C(_04554_),
    .Y(_04556_)
  );
  XOR2X1 _12392_ (
    .A(multiplier_0.reshi_10_ ),
    .B(_04555_),
    .Y(_04557_)
  );
  XNOR2X1 _12393_ (
    .A(_04502_),
    .B(_04503_),
    .Y(_04558_)
  );
  NAND2X1 _12394_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04558_),
    .Y(_04559_)
  );
  NAND2X1 _12395_ (
    .A(_04532_),
    .B(_04559_),
    .Y(_04560_)
  );
  NAND2X1 _12396_ (
    .A(_05068_),
    .B(_04560_),
    .Y(_04561_)
  );
  NAND3X1 _12397_ (
    .A(multiplier_0.reshi_9_ ),
    .B(_04532_),
    .C(_04559_),
    .Y(_04562_)
  );
  INVX1 _12398_ (
    .A(_04562_),
    .Y(_04563_)
  );
  XNOR2X1 _12399_ (
    .A(_05540_),
    .B(_04501_),
    .Y(_04564_)
  );
  OR2X1 _12400_ (
    .A(_05047_),
    .B(_04564_),
    .Y(_04565_)
  );
  OAI21X1 _12401_ (
    .A(_05047_),
    .B(_04564_),
    .C(_04532_),
    .Y(_04566_)
  );
  NAND3X1 _12402_ (
    .A(multiplier_0.reshi_8_ ),
    .B(_04532_),
    .C(_04565_),
    .Y(_04567_)
  );
  AOI21X1 _12403_ (
    .A(_04532_),
    .B(_04565_),
    .C(multiplier_0.reshi_8_ ),
    .Y(_04568_)
  );
  XOR2X1 _12404_ (
    .A(multiplier_0.reshi_8_ ),
    .B(_04566_),
    .Y(_04569_)
  );
  XNOR2X1 _12405_ (
    .A(_04499_),
    .B(_04500_),
    .Y(_04570_)
  );
  AND2X1 _12406_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04570_),
    .Y(_04571_)
  );
  NOR2X1 _12407_ (
    .A(_04531_),
    .B(_04571_),
    .Y(_04572_)
  );
  NOR3X1 _12408_ (
    .A(_05069_),
    .B(_04531_),
    .C(_04571_),
    .Y(_04573_)
  );
  NOR2X1 _12409_ (
    .A(multiplier_0.reshi_7_ ),
    .B(_04572_),
    .Y(_04574_)
  );
  OAI21X1 _12410_ (
    .A(_04531_),
    .B(_04571_),
    .C(_05069_),
    .Y(_04575_)
  );
  NOR2X1 _12411_ (
    .A(_04573_),
    .B(_04574_),
    .Y(_04576_)
  );
  XNOR2X1 _12412_ (
    .A(_05626_),
    .B(_04498_),
    .Y(_04577_)
  );
  MUX2X1 _12413_ (
    .A(_04529_),
    .B(_04577_),
    .S(_05047_),
    .Y(_04578_)
  );
  NAND2X1 _12414_ (
    .A(multiplier_0.reshi_6_ ),
    .B(_04578_),
    .Y(_04579_)
  );
  XNOR2X1 _12415_ (
    .A(multiplier_0.reshi_6_ ),
    .B(_04578_),
    .Y(_04580_)
  );
  XNOR2X1 _12416_ (
    .A(_05667_),
    .B(_04497_),
    .Y(_04581_)
  );
  MUX2X1 _12417_ (
    .A(_04536_),
    .B(_04581_),
    .S(_05047_),
    .Y(_04582_)
  );
  AND2X1 _12418_ (
    .A(multiplier_0.reshi_5_ ),
    .B(_04582_),
    .Y(_04583_)
  );
  NAND2X1 _12419_ (
    .A(multiplier_0.reshi_5_ ),
    .B(_04582_),
    .Y(_04584_)
  );
  XOR2X1 _12420_ (
    .A(_05713_),
    .B(_04496_),
    .Y(_04585_)
  );
  NAND2X1 _12421_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04585_),
    .Y(_04586_)
  );
  OAI21X1 _12422_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04542_),
    .C(_04586_),
    .Y(_04587_)
  );
  NAND2X1 _12423_ (
    .A(multiplier_0.reshi_4_ ),
    .B(_04587_),
    .Y(_04588_)
  );
  XNOR2X1 _12424_ (
    .A(multiplier_0.reshi_4_ ),
    .B(_04587_),
    .Y(_04589_)
  );
  XNOR2X1 _12425_ (
    .A(_05750_),
    .B(_04495_),
    .Y(_04590_)
  );
  MUX2X1 _12426_ (
    .A(_04547_),
    .B(_04590_),
    .S(_05047_),
    .Y(_04591_)
  );
  AND2X1 _12427_ (
    .A(multiplier_0.reshi_3_ ),
    .B(_04591_),
    .Y(_04592_)
  );
  NAND2X1 _12428_ (
    .A(multiplier_0.reshi_3_ ),
    .B(_04591_),
    .Y(_04593_)
  );
  OR2X1 _12429_ (
    .A(multiplier_0.reshi_3_ ),
    .B(_04591_),
    .Y(_04594_)
  );
  NAND2X1 _12430_ (
    .A(_04593_),
    .B(_04594_),
    .Y(_04595_)
  );
  XNOR2X1 _12431_ (
    .A(_05787_),
    .B(_04494_),
    .Y(_04596_)
  );
  MUX2X1 _12432_ (
    .A(_04553_),
    .B(_04596_),
    .S(_05047_),
    .Y(_04597_)
  );
  NAND2X1 _12433_ (
    .A(multiplier_0.reshi_2_ ),
    .B(_04597_),
    .Y(_04598_)
  );
  XNOR2X1 _12434_ (
    .A(multiplier_0.reshi_2_ ),
    .B(_04597_),
    .Y(_04599_)
  );
  XNOR2X1 _12435_ (
    .A(_04492_),
    .B(_04493_),
    .Y(_04600_)
  );
  MUX2X1 _12436_ (
    .A(_04558_),
    .B(_04600_),
    .S(_05047_),
    .Y(_04601_)
  );
  AND2X1 _12437_ (
    .A(multiplier_0.reshi_1_ ),
    .B(_04601_),
    .Y(_04602_)
  );
  NAND2X1 _12438_ (
    .A(multiplier_0.reshi_1_ ),
    .B(_04601_),
    .Y(_04603_)
  );
  OR2X1 _12439_ (
    .A(multiplier_0.reshi_1_ ),
    .B(_04601_),
    .Y(_04604_)
  );
  NAND2X1 _12440_ (
    .A(_04603_),
    .B(_04604_),
    .Y(_04605_)
  );
  XNOR2X1 _12441_ (
    .A(_04490_),
    .B(_04491_),
    .Y(_04606_)
  );
  NAND2X1 _12442_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04606_),
    .Y(_04607_)
  );
  OAI21X1 _12443_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04564_),
    .C(_04607_),
    .Y(_04608_)
  );
  NOR2X1 _12444_ (
    .A(_05070_),
    .B(_04608_),
    .Y(_04609_)
  );
  OR2X1 _12445_ (
    .A(_05070_),
    .B(_04608_),
    .Y(_04610_)
  );
  XNOR2X1 _12446_ (
    .A(_04488_),
    .B(_04489_),
    .Y(_04611_)
  );
  MUX2X1 _12447_ (
    .A(_04570_),
    .B(_04611_),
    .S(_05047_),
    .Y(_04612_)
  );
  AND2X1 _12448_ (
    .A(multiplier_0.reslo_15_ ),
    .B(_04612_),
    .Y(_04613_)
  );
  XOR2X1 _12449_ (
    .A(multiplier_0.reslo_15_ ),
    .B(_04612_),
    .Y(_04614_)
  );
  XOR2X1 _12450_ (
    .A(_04486_),
    .B(_04487_),
    .Y(_04615_)
  );
  NAND2X1 _12451_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04615_),
    .Y(_04616_)
  );
  OAI21X1 _12452_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04577_),
    .C(_04616_),
    .Y(_04617_)
  );
  NAND2X1 _12453_ (
    .A(multiplier_0.reslo_14_ ),
    .B(_04617_),
    .Y(_04618_)
  );
  XNOR2X1 _12454_ (
    .A(multiplier_0.reslo_14_ ),
    .B(_04617_),
    .Y(_04619_)
  );
  XNOR2X1 _12455_ (
    .A(_04483_),
    .B(_04485_),
    .Y(_04620_)
  );
  NAND2X1 _12456_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04620_),
    .Y(_04621_)
  );
  OAI21X1 _12457_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04581_),
    .C(_04621_),
    .Y(_04622_)
  );
  AND2X1 _12458_ (
    .A(multiplier_0.reslo_13_ ),
    .B(_04622_),
    .Y(_04623_)
  );
  XOR2X1 _12459_ (
    .A(multiplier_0.reslo_13_ ),
    .B(_04622_),
    .Y(_04624_)
  );
  XOR2X1 _12460_ (
    .A(_04480_),
    .B(_04482_),
    .Y(_04625_)
  );
  NAND2X1 _12461_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04625_),
    .Y(_04626_)
  );
  OAI21X1 _12462_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04585_),
    .C(_04626_),
    .Y(_04627_)
  );
  NOR2X1 _12463_ (
    .A(_05071_),
    .B(_04627_),
    .Y(_04628_)
  );
  OR2X1 _12464_ (
    .A(_05071_),
    .B(_04627_),
    .Y(_04629_)
  );
  AND2X1 _12465_ (
    .A(_05071_),
    .B(_04627_),
    .Y(_04630_)
  );
  NOR2X1 _12466_ (
    .A(_04628_),
    .B(_04630_),
    .Y(_04631_)
  );
  XNOR2X1 _12467_ (
    .A(_04477_),
    .B(_04479_),
    .Y(_04632_)
  );
  NAND2X1 _12468_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04632_),
    .Y(_04633_)
  );
  OAI21X1 _12469_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04590_),
    .C(_04633_),
    .Y(_04634_)
  );
  AND2X1 _12470_ (
    .A(multiplier_0.reslo_11_ ),
    .B(_04634_),
    .Y(_04635_)
  );
  NAND2X1 _12471_ (
    .A(_04474_),
    .B(_04476_),
    .Y(_04636_)
  );
  NAND2X1 _12472_ (
    .A(_04478_),
    .B(_04636_),
    .Y(_04637_)
  );
  MUX2X1 _12473_ (
    .A(_04596_),
    .B(_04637_),
    .S(_05047_),
    .Y(_04638_)
  );
  NAND2X1 _12474_ (
    .A(multiplier_0.reslo_10_ ),
    .B(_04638_),
    .Y(_04639_)
  );
  XNOR2X1 _12475_ (
    .A(multiplier_0.reslo_10_ ),
    .B(_04638_),
    .Y(_04640_)
  );
  AOI22X1 _12476_ (
    .A(multiplier_0.op1_0_ ),
    .B(_05159_),
    .C(_05169_),
    .D(multiplier_0.op1_1_ ),
    .Y(_04641_)
  );
  NOR2X1 _12477_ (
    .A(_04475_),
    .B(_04641_),
    .Y(_04642_)
  );
  NAND2X1 _12478_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04642_),
    .Y(_04643_)
  );
  OAI21X1 _12479_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04600_),
    .C(_04643_),
    .Y(_04644_)
  );
  AND2X1 _12480_ (
    .A(multiplier_0.reslo_9_ ),
    .B(_04644_),
    .Y(_04645_)
  );
  AOI21X1 _12481_ (
    .A(multiplier_0.op2_8_ ),
    .B(multiplier_0.op1_0_ ),
    .C(_05047_),
    .Y(_04646_)
  );
  AOI21X1 _12482_ (
    .A(_05047_),
    .B(_04606_),
    .C(_04646_),
    .Y(_04647_)
  );
  NAND2X1 _12483_ (
    .A(multiplier_0.reslo_8_ ),
    .B(_04647_),
    .Y(_04648_)
  );
  NOR2X1 _12484_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04611_),
    .Y(_04649_)
  );
  AND2X1 _12485_ (
    .A(multiplier_0.reslo_7_ ),
    .B(_04649_),
    .Y(_04650_)
  );
  XOR2X1 _12486_ (
    .A(multiplier_0.reslo_7_ ),
    .B(_04649_),
    .Y(_04651_)
  );
  NAND2X1 _12487_ (
    .A(_05047_),
    .B(_04615_),
    .Y(_04652_)
  );
  NAND3X1 _12488_ (
    .A(_05047_),
    .B(multiplier_0.reslo_6_ ),
    .C(_04615_),
    .Y(_04653_)
  );
  AOI21X1 _12489_ (
    .A(_05047_),
    .B(_04615_),
    .C(multiplier_0.reslo_6_ ),
    .Y(_04654_)
  );
  XNOR2X1 _12490_ (
    .A(multiplier_0.reslo_6_ ),
    .B(_04652_),
    .Y(_04655_)
  );
  NAND2X1 _12491_ (
    .A(_05047_),
    .B(_04620_),
    .Y(_04656_)
  );
  NOR2X1 _12492_ (
    .A(_05072_),
    .B(_04656_),
    .Y(_04657_)
  );
  XNOR2X1 _12493_ (
    .A(multiplier_0.reslo_5_ ),
    .B(_04656_),
    .Y(_04658_)
  );
  NOR2X1 _12494_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04625_),
    .Y(_04659_)
  );
  NAND2X1 _12495_ (
    .A(multiplier_0.reslo_4_ ),
    .B(_04659_),
    .Y(_04660_)
  );
  XNOR2X1 _12496_ (
    .A(multiplier_0.reslo_4_ ),
    .B(_04659_),
    .Y(_04661_)
  );
  NAND3X1 _12497_ (
    .A(_05047_),
    .B(multiplier_0.reslo_3_ ),
    .C(_04632_),
    .Y(_04662_)
  );
  INVX1 _12498_ (
    .A(_04662_),
    .Y(_04663_)
  );
  AOI21X1 _12499_ (
    .A(_05047_),
    .B(_04632_),
    .C(multiplier_0.reslo_3_ ),
    .Y(_04664_)
  );
  NOR2X1 _12500_ (
    .A(_04663_),
    .B(_04664_),
    .Y(_04665_)
  );
  NOR2X1 _12501_ (
    .A(multiplier_0.cycle_0_ ),
    .B(_04637_),
    .Y(_04666_)
  );
  NAND2X1 _12502_ (
    .A(multiplier_0.reslo_2_ ),
    .B(_04666_),
    .Y(_04667_)
  );
  AND2X1 _12503_ (
    .A(_05047_),
    .B(_04642_),
    .Y(_04668_)
  );
  NAND2X1 _12504_ (
    .A(multiplier_0.reslo_1_ ),
    .B(_04668_),
    .Y(_04669_)
  );
  NAND2X1 _12505_ (
    .A(multiplier_0.reslo_0_ ),
    .B(_04473_),
    .Y(_04670_)
  );
  XNOR2X1 _12506_ (
    .A(multiplier_0.reslo_1_ ),
    .B(_04668_),
    .Y(_04671_)
  );
  OAI21X1 _12507_ (
    .A(_04670_),
    .B(_04671_),
    .C(_04669_),
    .Y(_04672_)
  );
  XOR2X1 _12508_ (
    .A(multiplier_0.reslo_2_ ),
    .B(_04666_),
    .Y(_04673_)
  );
  NAND2X1 _12509_ (
    .A(_04672_),
    .B(_04673_),
    .Y(_04674_)
  );
  NAND2X1 _12510_ (
    .A(_04667_),
    .B(_04674_),
    .Y(_04675_)
  );
  AOI21X1 _12511_ (
    .A(_04665_),
    .B(_04675_),
    .C(_04663_),
    .Y(_04676_)
  );
  OAI21X1 _12512_ (
    .A(_04661_),
    .B(_04676_),
    .C(_04660_),
    .Y(_04677_)
  );
  AOI21X1 _12513_ (
    .A(_04658_),
    .B(_04677_),
    .C(_04657_),
    .Y(_04678_)
  );
  OAI21X1 _12514_ (
    .A(_04654_),
    .B(_04678_),
    .C(_04653_),
    .Y(_04679_)
  );
  AOI21X1 _12515_ (
    .A(_04651_),
    .B(_04679_),
    .C(_04650_),
    .Y(_04680_)
  );
  XNOR2X1 _12516_ (
    .A(multiplier_0.reslo_8_ ),
    .B(_04647_),
    .Y(_04681_)
  );
  OAI21X1 _12517_ (
    .A(_04680_),
    .B(_04681_),
    .C(_04648_),
    .Y(_04682_)
  );
  XOR2X1 _12518_ (
    .A(multiplier_0.reslo_9_ ),
    .B(_04644_),
    .Y(_04683_)
  );
  AOI21X1 _12519_ (
    .A(_04682_),
    .B(_04683_),
    .C(_04645_),
    .Y(_04684_)
  );
  OAI21X1 _12520_ (
    .A(_04640_),
    .B(_04684_),
    .C(_04639_),
    .Y(_04685_)
  );
  XOR2X1 _12521_ (
    .A(multiplier_0.reslo_11_ ),
    .B(_04634_),
    .Y(_04686_)
  );
  AOI21X1 _12522_ (
    .A(_04685_),
    .B(_04686_),
    .C(_04635_),
    .Y(_04687_)
  );
  OAI21X1 _12523_ (
    .A(_04630_),
    .B(_04687_),
    .C(_04629_),
    .Y(_04688_)
  );
  AOI21X1 _12524_ (
    .A(_04624_),
    .B(_04688_),
    .C(_04623_),
    .Y(_04689_)
  );
  OAI21X1 _12525_ (
    .A(_04619_),
    .B(_04689_),
    .C(_04618_),
    .Y(_04690_)
  );
  AOI21X1 _12526_ (
    .A(_04614_),
    .B(_04690_),
    .C(_04613_),
    .Y(_04691_)
  );
  AND2X1 _12527_ (
    .A(_05070_),
    .B(_04608_),
    .Y(_04692_)
  );
  NOR2X1 _12528_ (
    .A(_04609_),
    .B(_04692_),
    .Y(_04693_)
  );
  OAI21X1 _12529_ (
    .A(_04691_),
    .B(_04692_),
    .C(_04610_),
    .Y(_04694_)
  );
  AOI21X1 _12530_ (
    .A(_04604_),
    .B(_04694_),
    .C(_04602_),
    .Y(_04695_)
  );
  OAI21X1 _12531_ (
    .A(_04599_),
    .B(_04695_),
    .C(_04598_),
    .Y(_04696_)
  );
  AOI21X1 _12532_ (
    .A(_04594_),
    .B(_04696_),
    .C(_04592_),
    .Y(_04697_)
  );
  OAI21X1 _12533_ (
    .A(_04589_),
    .B(_04697_),
    .C(_04588_),
    .Y(_04698_)
  );
  OR2X1 _12534_ (
    .A(multiplier_0.reshi_5_ ),
    .B(_04582_),
    .Y(_04699_)
  );
  NAND2X1 _12535_ (
    .A(_04584_),
    .B(_04699_),
    .Y(_04700_)
  );
  AOI21X1 _12536_ (
    .A(_04698_),
    .B(_04699_),
    .C(_04583_),
    .Y(_04701_)
  );
  OAI21X1 _12537_ (
    .A(_04580_),
    .B(_04701_),
    .C(_04579_),
    .Y(_04702_)
  );
  AOI21X1 _12538_ (
    .A(_04575_),
    .B(_04702_),
    .C(_04573_),
    .Y(_04703_)
  );
  OAI21X1 _12539_ (
    .A(_04568_),
    .B(_04703_),
    .C(_04567_),
    .Y(_04704_)
  );
  AOI21X1 _12540_ (
    .A(_04561_),
    .B(_04704_),
    .C(_04563_),
    .Y(_04705_)
  );
  OAI21X1 _12541_ (
    .A(_04557_),
    .B(_04705_),
    .C(_04556_),
    .Y(_04706_)
  );
  AOI21X1 _12542_ (
    .A(_04550_),
    .B(_04706_),
    .C(_04552_),
    .Y(_04707_)
  );
  OAI21X1 _12543_ (
    .A(_04546_),
    .B(_04707_),
    .C(_04545_),
    .Y(_04708_)
  );
  OAI21X1 _12544_ (
    .A(_04540_),
    .B(_04708_),
    .C(_04541_),
    .Y(_04709_)
  );
  OAI21X1 _12545_ (
    .A(_04535_),
    .B(_04709_),
    .C(_04534_),
    .Y(_04710_)
  );
  NAND2X1 _12546_ (
    .A(_04528_),
    .B(_04710_),
    .Y(_04711_)
  );
  XNOR2X1 _12547_ (
    .A(_04528_),
    .B(_04710_),
    .Y(_04712_)
  );
  NOR2X1 _12548_ (
    .A(_05049_),
    .B(_04712_),
    .Y(_04713_)
  );
  AOI21X1 _12549_ (
    .A(multiplier_0.reshi_15_ ),
    .B(_04526_),
    .C(multiplier_0.sumext_0_ ),
    .Y(_04714_)
  );
  AOI21X1 _12550_ (
    .A(_04711_),
    .B(_04714_),
    .C(multiplier_0.sign_sel ),
    .Y(_04715_)
  );
  NOR2X1 _12551_ (
    .A(_04713_),
    .B(_04715_),
    .Y(_04716_)
  );
  NOR2X1 _12552_ (
    .A(_05045_),
    .B(_00109_),
    .Y(_04717_)
  );
  NAND3X1 _12553_ (
    .A(_00103_),
    .B(_05044_),
    .C(_04717_),
    .Y(_04718_)
  );
  NOR2X1 _12554_ (
    .A(_00108_),
    .B(_00098_),
    .Y(_04719_)
  );
  NOR2X1 _12555_ (
    .A(_05043_),
    .B(_00105_),
    .Y(_04720_)
  );
  NAND3X1 _12556_ (
    .A(_05083_),
    .B(_04719_),
    .C(_04720_),
    .Y(_04721_)
  );
  NOR2X1 _12557_ (
    .A(_04718_),
    .B(_04721_),
    .Y(_04722_)
  );
  OAI21X1 _12558_ (
    .A(_00127_),
    .B(_00128_),
    .C(_04722_),
    .Y(_04723_)
  );
  OR2X1 _12559_ (
    .A(_05080_),
    .B(_04723_),
    .Y(_04724_)
  );
  NOR2X1 _12560_ (
    .A(_00106_),
    .B(_05081_),
    .Y(_04725_)
  );
  NOR2X1 _12561_ (
    .A(_00105_),
    .B(_00098_),
    .Y(_04726_)
  );
  NAND3X1 _12562_ (
    .A(_00104_),
    .B(_04725_),
    .C(_04726_),
    .Y(_04727_)
  );
  NAND2X1 _12563_ (
    .A(_00103_),
    .B(_00107_),
    .Y(_04728_)
  );
  NOR2X1 _12564_ (
    .A(_00109_),
    .B(_04728_),
    .Y(_04729_)
  );
  NOR2X1 _12565_ (
    .A(_00108_),
    .B(_05082_),
    .Y(_04730_)
  );
  NAND2X1 _12566_ (
    .A(_04729_),
    .B(_04730_),
    .Y(_04731_)
  );
  NOR2X1 _12567_ (
    .A(_04727_),
    .B(_04731_),
    .Y(_04732_)
  );
  OAI21X1 _12568_ (
    .A(_00127_),
    .B(_00128_),
    .C(_04732_),
    .Y(_04733_)
  );
  OR2X1 _12569_ (
    .A(_05080_),
    .B(_04733_),
    .Y(_04734_)
  );
  OAI21X1 _12570_ (
    .A(multiplier_0.sumext_0_ ),
    .B(_05095_),
    .C(_04724_),
    .Y(_04735_)
  );
  AOI21X1 _12571_ (
    .A(_05095_),
    .B(_04716_),
    .C(_04735_),
    .Y(_04439_)
  );
  NOR2X1 _12572_ (
    .A(_05094_),
    .B(_04713_),
    .Y(_04736_)
  );
  OAI21X1 _12573_ (
    .A(multiplier_0.sumext_10_ ),
    .B(_05095_),
    .C(_05093_),
    .Y(_04737_)
  );
  NOR2X1 _12574_ (
    .A(_04736_),
    .B(_04737_),
    .Y(_04440_)
  );
  OAI21X1 _12575_ (
    .A(_05080_),
    .B(_04733_),
    .C(_05058_),
    .Y(_04738_)
  );
  OAI21X1 _12576_ (
    .A(_00110_),
    .B(_04734_),
    .C(_04738_),
    .Y(_04739_)
  );
  INVX1 _12577_ (
    .A(_04739_),
    .Y(_04390_)
  );
  OAI21X1 _12578_ (
    .A(_05080_),
    .B(_04733_),
    .C(_05057_),
    .Y(_04740_)
  );
  OAI21X1 _12579_ (
    .A(_00117_),
    .B(_04734_),
    .C(_04740_),
    .Y(_04741_)
  );
  INVX1 _12580_ (
    .A(_04741_),
    .Y(_04397_)
  );
  OAI21X1 _12581_ (
    .A(_05080_),
    .B(_04733_),
    .C(_05056_),
    .Y(_04742_)
  );
  OAI21X1 _12582_ (
    .A(_00118_),
    .B(_04734_),
    .C(_04742_),
    .Y(_04743_)
  );
  INVX1 _12583_ (
    .A(_04743_),
    .Y(_04398_)
  );
  OAI21X1 _12584_ (
    .A(_05080_),
    .B(_04733_),
    .C(_05055_),
    .Y(_04744_)
  );
  OAI21X1 _12585_ (
    .A(_00119_),
    .B(_04734_),
    .C(_04744_),
    .Y(_04745_)
  );
  INVX1 _12586_ (
    .A(_04745_),
    .Y(_04399_)
  );
  OAI21X1 _12587_ (
    .A(_05080_),
    .B(_04733_),
    .C(_05054_),
    .Y(_04746_)
  );
  OAI21X1 _12588_ (
    .A(_00120_),
    .B(_04734_),
    .C(_04746_),
    .Y(_04747_)
  );
  INVX1 _12589_ (
    .A(_04747_),
    .Y(_04400_)
  );
  OAI21X1 _12590_ (
    .A(_05080_),
    .B(_04733_),
    .C(_05053_),
    .Y(_04748_)
  );
  OAI21X1 _12591_ (
    .A(_00121_),
    .B(_04734_),
    .C(_04748_),
    .Y(_04749_)
  );
  INVX1 _12592_ (
    .A(_04749_),
    .Y(_04401_)
  );
  OAI21X1 _12593_ (
    .A(_05080_),
    .B(_04733_),
    .C(_05052_),
    .Y(_04750_)
  );
  OAI21X1 _12594_ (
    .A(_00122_),
    .B(_04734_),
    .C(_04750_),
    .Y(_04751_)
  );
  INVX1 _12595_ (
    .A(_04751_),
    .Y(_04402_)
  );
  OAI21X1 _12596_ (
    .A(_05080_),
    .B(_04733_),
    .C(_05051_),
    .Y(_04752_)
  );
  OAI21X1 _12597_ (
    .A(_00123_),
    .B(_04734_),
    .C(_04752_),
    .Y(_04753_)
  );
  INVX1 _12598_ (
    .A(_04753_),
    .Y(_04403_)
  );
  OAI21X1 _12599_ (
    .A(_05080_),
    .B(_05092_),
    .C(multiplier_0.op2_8_ ),
    .Y(_04754_)
  );
  NAND2X1 _12600_ (
    .A(_00128_),
    .B(_00124_),
    .Y(_04755_)
  );
  OAI21X1 _12601_ (
    .A(_04724_),
    .B(_04755_),
    .C(_04754_),
    .Y(_04404_)
  );
  OAI21X1 _12602_ (
    .A(_05080_),
    .B(_05092_),
    .C(multiplier_0.op2_9_ ),
    .Y(_04756_)
  );
  NAND2X1 _12603_ (
    .A(_00128_),
    .B(_00125_),
    .Y(_04757_)
  );
  OAI21X1 _12604_ (
    .A(_04724_),
    .B(_04757_),
    .C(_04756_),
    .Y(_04405_)
  );
  OAI21X1 _12605_ (
    .A(_05080_),
    .B(_05092_),
    .C(multiplier_0.op2_10_ ),
    .Y(_04758_)
  );
  NAND2X1 _12606_ (
    .A(_00128_),
    .B(_00111_),
    .Y(_04759_)
  );
  OAI21X1 _12607_ (
    .A(_04724_),
    .B(_04759_),
    .C(_04758_),
    .Y(_04391_)
  );
  OAI21X1 _12608_ (
    .A(_05080_),
    .B(_05092_),
    .C(multiplier_0.op2_11_ ),
    .Y(_04760_)
  );
  NAND2X1 _12609_ (
    .A(_00128_),
    .B(_00112_),
    .Y(_04761_)
  );
  OAI21X1 _12610_ (
    .A(_04724_),
    .B(_04761_),
    .C(_04760_),
    .Y(_04392_)
  );
  OAI21X1 _12611_ (
    .A(_05080_),
    .B(_05092_),
    .C(multiplier_0.op2_12_ ),
    .Y(_04762_)
  );
  NAND2X1 _12612_ (
    .A(_00128_),
    .B(_00113_),
    .Y(_04763_)
  );
  OAI21X1 _12613_ (
    .A(_04724_),
    .B(_04763_),
    .C(_04762_),
    .Y(_04393_)
  );
  OAI21X1 _12614_ (
    .A(_05080_),
    .B(_05092_),
    .C(multiplier_0.op2_13_ ),
    .Y(_04764_)
  );
  NAND2X1 _12615_ (
    .A(_00128_),
    .B(_00114_),
    .Y(_04765_)
  );
  OAI21X1 _12616_ (
    .A(_04724_),
    .B(_04765_),
    .C(_04764_),
    .Y(_04394_)
  );
  OAI21X1 _12617_ (
    .A(_05080_),
    .B(_05092_),
    .C(multiplier_0.op2_14_ ),
    .Y(_04766_)
  );
  NAND2X1 _12618_ (
    .A(_00128_),
    .B(_00115_),
    .Y(_04767_)
  );
  OAI21X1 _12619_ (
    .A(_04724_),
    .B(_04767_),
    .C(_04766_),
    .Y(_04395_)
  );
  OAI21X1 _12620_ (
    .A(_05080_),
    .B(_05092_),
    .C(multiplier_0.op2_15_ ),
    .Y(_04768_)
  );
  NAND2X1 _12621_ (
    .A(_00128_),
    .B(_00116_),
    .Y(_04769_)
  );
  OAI21X1 _12622_ (
    .A(_04724_),
    .B(_04769_),
    .C(_04768_),
    .Y(_04396_)
  );
  NAND2X1 _12623_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04473_),
    .Y(_04770_)
  );
  XNOR2X1 _12624_ (
    .A(multiplier_0.reslo_0_ ),
    .B(_04770_),
    .Y(_04771_)
  );
  NAND2X1 _12625_ (
    .A(_00097_),
    .B(_00102_),
    .Y(_04772_)
  );
  OR2X1 _12626_ (
    .A(_00101_),
    .B(_04772_),
    .Y(_04773_)
  );
  OR2X1 _12627_ (
    .A(_05092_),
    .B(_04773_),
    .Y(_04774_)
  );
  INVX1 _12628_ (
    .A(_04774_),
    .Y(_04775_)
  );
  NOR2X1 _12629_ (
    .A(multiplier_0.acc_sel ),
    .B(_04734_),
    .Y(_04776_)
  );
  NOR2X1 _12630_ (
    .A(_04733_),
    .B(_04773_),
    .Y(_04777_)
  );
  NOR2X1 _12631_ (
    .A(_04776_),
    .B(_04777_),
    .Y(_04778_)
  );
  INVX1 _12632_ (
    .A(_04778_),
    .Y(_04779_)
  );
  NAND2X1 _12633_ (
    .A(_04771_),
    .B(_04778_),
    .Y(_04780_)
  );
  OAI21X1 _12634_ (
    .A(_05073_),
    .B(_04774_),
    .C(_04780_),
    .Y(_04422_)
  );
  XNOR2X1 _12635_ (
    .A(_04670_),
    .B(_04671_),
    .Y(_04781_)
  );
  NAND2X1 _12636_ (
    .A(multiplier_0.reslo_1_ ),
    .B(_05094_),
    .Y(_04782_)
  );
  OAI21X1 _12637_ (
    .A(_05094_),
    .B(_04781_),
    .C(_04782_),
    .Y(_04783_)
  );
  NAND2X1 _12638_ (
    .A(_04778_),
    .B(_04783_),
    .Y(_04784_)
  );
  OAI21X1 _12639_ (
    .A(_05074_),
    .B(_04774_),
    .C(_04784_),
    .Y(_04429_)
  );
  XNOR2X1 _12640_ (
    .A(_04672_),
    .B(_04673_),
    .Y(_04785_)
  );
  NAND2X1 _12641_ (
    .A(multiplier_0.reslo_2_ ),
    .B(_05094_),
    .Y(_04786_)
  );
  OAI21X1 _12642_ (
    .A(_05094_),
    .B(_04785_),
    .C(_04786_),
    .Y(_04787_)
  );
  NAND2X1 _12643_ (
    .A(_04778_),
    .B(_04787_),
    .Y(_04788_)
  );
  OAI21X1 _12644_ (
    .A(_05075_),
    .B(_04774_),
    .C(_04788_),
    .Y(_04430_)
  );
  XNOR2X1 _12645_ (
    .A(_04665_),
    .B(_04675_),
    .Y(_04789_)
  );
  NAND2X1 _12646_ (
    .A(multiplier_0.reslo_3_ ),
    .B(_05094_),
    .Y(_04790_)
  );
  OAI21X1 _12647_ (
    .A(_05094_),
    .B(_04789_),
    .C(_04790_),
    .Y(_04791_)
  );
  NAND2X1 _12648_ (
    .A(_04778_),
    .B(_04791_),
    .Y(_04792_)
  );
  OAI21X1 _12649_ (
    .A(_05076_),
    .B(_04774_),
    .C(_04792_),
    .Y(_04431_)
  );
  XNOR2X1 _12650_ (
    .A(_04661_),
    .B(_04676_),
    .Y(_04793_)
  );
  OAI21X1 _12651_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_04793_),
    .Y(_04794_)
  );
  OAI21X1 _12652_ (
    .A(multiplier_0.reslo_4_ ),
    .B(_05095_),
    .C(_04794_),
    .Y(_04795_)
  );
  NAND2X1 _12653_ (
    .A(_00120_),
    .B(_04775_),
    .Y(_04796_)
  );
  OAI21X1 _12654_ (
    .A(_04779_),
    .B(_04795_),
    .C(_04796_),
    .Y(_04432_)
  );
  XNOR2X1 _12655_ (
    .A(_04658_),
    .B(_04677_),
    .Y(_04797_)
  );
  OAI21X1 _12656_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_04797_),
    .Y(_04798_)
  );
  OAI21X1 _12657_ (
    .A(multiplier_0.reslo_5_ ),
    .B(_05095_),
    .C(_04798_),
    .Y(_04799_)
  );
  NAND2X1 _12658_ (
    .A(_00121_),
    .B(_04775_),
    .Y(_04800_)
  );
  OAI21X1 _12659_ (
    .A(_04779_),
    .B(_04799_),
    .C(_04800_),
    .Y(_04433_)
  );
  XOR2X1 _12660_ (
    .A(_04655_),
    .B(_04678_),
    .Y(_04801_)
  );
  NAND2X1 _12661_ (
    .A(multiplier_0.reslo_6_ ),
    .B(_05094_),
    .Y(_04802_)
  );
  OAI21X1 _12662_ (
    .A(_05094_),
    .B(_04801_),
    .C(_04802_),
    .Y(_04803_)
  );
  NAND2X1 _12663_ (
    .A(_04778_),
    .B(_04803_),
    .Y(_04804_)
  );
  OAI21X1 _12664_ (
    .A(_05077_),
    .B(_04774_),
    .C(_04804_),
    .Y(_04434_)
  );
  XNOR2X1 _12665_ (
    .A(_04651_),
    .B(_04679_),
    .Y(_04805_)
  );
  OAI21X1 _12666_ (
    .A(multiplier_0.cycle_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_04805_),
    .Y(_04806_)
  );
  OAI21X1 _12667_ (
    .A(multiplier_0.reslo_7_ ),
    .B(_05095_),
    .C(_04806_),
    .Y(_04807_)
  );
  NAND2X1 _12668_ (
    .A(_00123_),
    .B(_04775_),
    .Y(_04808_)
  );
  OAI21X1 _12669_ (
    .A(_04779_),
    .B(_04807_),
    .C(_04808_),
    .Y(_04435_)
  );
  XNOR2X1 _12670_ (
    .A(_04680_),
    .B(_04681_),
    .Y(_04809_)
  );
  AOI21X1 _12671_ (
    .A(_05095_),
    .B(_04809_),
    .C(_04779_),
    .Y(_04810_)
  );
  OAI21X1 _12672_ (
    .A(multiplier_0.reslo_8_ ),
    .B(_05095_),
    .C(_04810_),
    .Y(_04811_)
  );
  OAI21X1 _12673_ (
    .A(_04755_),
    .B(_04774_),
    .C(_04811_),
    .Y(_04436_)
  );
  XNOR2X1 _12674_ (
    .A(_04682_),
    .B(_04683_),
    .Y(_04812_)
  );
  OAI21X1 _12675_ (
    .A(multiplier_0.reslo_9_ ),
    .B(_05095_),
    .C(_04778_),
    .Y(_04813_)
  );
  AOI21X1 _12676_ (
    .A(_05095_),
    .B(_04812_),
    .C(_04813_),
    .Y(_04814_)
  );
  INVX1 _12677_ (
    .A(_04814_),
    .Y(_04815_)
  );
  OAI21X1 _12678_ (
    .A(_04757_),
    .B(_04774_),
    .C(_04815_),
    .Y(_04437_)
  );
  XNOR2X1 _12679_ (
    .A(_04640_),
    .B(_04684_),
    .Y(_04816_)
  );
  AOI21X1 _12680_ (
    .A(_05095_),
    .B(_04816_),
    .C(_04779_),
    .Y(_04817_)
  );
  OAI21X1 _12681_ (
    .A(multiplier_0.reslo_10_ ),
    .B(_05095_),
    .C(_04817_),
    .Y(_04818_)
  );
  OAI21X1 _12682_ (
    .A(_04759_),
    .B(_04774_),
    .C(_04818_),
    .Y(_04423_)
  );
  XNOR2X1 _12683_ (
    .A(_04685_),
    .B(_04686_),
    .Y(_04819_)
  );
  AOI21X1 _12684_ (
    .A(_05095_),
    .B(_04819_),
    .C(_04779_),
    .Y(_04820_)
  );
  OAI21X1 _12685_ (
    .A(multiplier_0.reslo_11_ ),
    .B(_05095_),
    .C(_04820_),
    .Y(_04821_)
  );
  OAI21X1 _12686_ (
    .A(_04761_),
    .B(_04774_),
    .C(_04821_),
    .Y(_04424_)
  );
  XOR2X1 _12687_ (
    .A(_04631_),
    .B(_04687_),
    .Y(_04822_)
  );
  OAI21X1 _12688_ (
    .A(multiplier_0.reslo_12_ ),
    .B(_05095_),
    .C(_04778_),
    .Y(_04823_)
  );
  AOI21X1 _12689_ (
    .A(_05095_),
    .B(_04822_),
    .C(_04823_),
    .Y(_04824_)
  );
  INVX1 _12690_ (
    .A(_04824_),
    .Y(_04825_)
  );
  OAI21X1 _12691_ (
    .A(_04763_),
    .B(_04774_),
    .C(_04825_),
    .Y(_04425_)
  );
  XNOR2X1 _12692_ (
    .A(_04624_),
    .B(_04688_),
    .Y(_04826_)
  );
  OAI21X1 _12693_ (
    .A(multiplier_0.reslo_13_ ),
    .B(_05095_),
    .C(_04778_),
    .Y(_04827_)
  );
  AOI21X1 _12694_ (
    .A(_05095_),
    .B(_04826_),
    .C(_04827_),
    .Y(_04828_)
  );
  INVX1 _12695_ (
    .A(_04828_),
    .Y(_04829_)
  );
  OAI21X1 _12696_ (
    .A(_04765_),
    .B(_04774_),
    .C(_04829_),
    .Y(_04426_)
  );
  XNOR2X1 _12697_ (
    .A(_04619_),
    .B(_04689_),
    .Y(_04830_)
  );
  AOI21X1 _12698_ (
    .A(_05095_),
    .B(_04830_),
    .C(_04779_),
    .Y(_04831_)
  );
  OAI21X1 _12699_ (
    .A(multiplier_0.reslo_14_ ),
    .B(_05095_),
    .C(_04831_),
    .Y(_04832_)
  );
  OAI21X1 _12700_ (
    .A(_04767_),
    .B(_04774_),
    .C(_04832_),
    .Y(_04427_)
  );
  XNOR2X1 _12701_ (
    .A(_04614_),
    .B(_04690_),
    .Y(_04833_)
  );
  OAI21X1 _12702_ (
    .A(multiplier_0.reslo_15_ ),
    .B(_05095_),
    .C(_04778_),
    .Y(_04834_)
  );
  AOI21X1 _12703_ (
    .A(_05095_),
    .B(_04833_),
    .C(_04834_),
    .Y(_04835_)
  );
  INVX1 _12704_ (
    .A(_04835_),
    .Y(_04836_)
  );
  OAI21X1 _12705_ (
    .A(_04769_),
    .B(_04774_),
    .C(_04836_),
    .Y(_04428_)
  );
  XOR2X1 _12706_ (
    .A(_04691_),
    .B(_04693_),
    .Y(_04837_)
  );
  NAND3X1 _12707_ (
    .A(_00101_),
    .B(_05042_),
    .C(_00102_),
    .Y(_04838_)
  );
  NOR2X1 _12708_ (
    .A(_05092_),
    .B(_04838_),
    .Y(_04839_)
  );
  NOR2X1 _12709_ (
    .A(_04733_),
    .B(_04838_),
    .Y(_04840_)
  );
  NOR2X1 _12710_ (
    .A(_04776_),
    .B(_04840_),
    .Y(_04841_)
  );
  OR2X1 _12711_ (
    .A(_04723_),
    .B(_04838_),
    .Y(_04842_)
  );
  OAI21X1 _12712_ (
    .A(multiplier_0.acc_sel ),
    .B(_04724_),
    .C(_04842_),
    .Y(_04843_)
  );
  AOI21X1 _12713_ (
    .A(_05095_),
    .B(_04837_),
    .C(_04843_),
    .Y(_04844_)
  );
  OAI21X1 _12714_ (
    .A(multiplier_0.reshi_0_ ),
    .B(_05095_),
    .C(_04844_),
    .Y(_04845_)
  );
  OAI21X1 _12715_ (
    .A(_05073_),
    .B(_04842_),
    .C(_04845_),
    .Y(_04406_)
  );
  XOR2X1 _12716_ (
    .A(_04605_),
    .B(_04694_),
    .Y(_04846_)
  );
  OAI21X1 _12717_ (
    .A(multiplier_0.reshi_1_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04847_)
  );
  AOI21X1 _12718_ (
    .A(_05095_),
    .B(_04846_),
    .C(_04847_),
    .Y(_04848_)
  );
  AOI21X1 _12719_ (
    .A(_00117_),
    .B(_04839_),
    .C(_04848_),
    .Y(_04849_)
  );
  INVX1 _12720_ (
    .A(_04849_),
    .Y(_04413_)
  );
  XNOR2X1 _12721_ (
    .A(_04599_),
    .B(_04695_),
    .Y(_04850_)
  );
  OAI21X1 _12722_ (
    .A(multiplier_0.reshi_2_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04851_)
  );
  AOI21X1 _12723_ (
    .A(_05095_),
    .B(_04850_),
    .C(_04851_),
    .Y(_04852_)
  );
  AOI21X1 _12724_ (
    .A(_00118_),
    .B(_04839_),
    .C(_04852_),
    .Y(_04853_)
  );
  INVX1 _12725_ (
    .A(_04853_),
    .Y(_04414_)
  );
  XOR2X1 _12726_ (
    .A(_04595_),
    .B(_04696_),
    .Y(_04854_)
  );
  OAI21X1 _12727_ (
    .A(multiplier_0.reshi_3_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04855_)
  );
  AOI21X1 _12728_ (
    .A(_05095_),
    .B(_04854_),
    .C(_04855_),
    .Y(_04856_)
  );
  AOI21X1 _12729_ (
    .A(_00119_),
    .B(_04839_),
    .C(_04856_),
    .Y(_04857_)
  );
  INVX1 _12730_ (
    .A(_04857_),
    .Y(_04415_)
  );
  XNOR2X1 _12731_ (
    .A(_04589_),
    .B(_04697_),
    .Y(_04858_)
  );
  OAI21X1 _12732_ (
    .A(multiplier_0.reshi_4_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04859_)
  );
  AOI21X1 _12733_ (
    .A(_05095_),
    .B(_04858_),
    .C(_04859_),
    .Y(_04860_)
  );
  AOI21X1 _12734_ (
    .A(_00120_),
    .B(_04839_),
    .C(_04860_),
    .Y(_04861_)
  );
  INVX1 _12735_ (
    .A(_04861_),
    .Y(_04416_)
  );
  XNOR2X1 _12736_ (
    .A(_04698_),
    .B(_04700_),
    .Y(_04862_)
  );
  NOR2X1 _12737_ (
    .A(_05094_),
    .B(_04862_),
    .Y(_04863_)
  );
  OAI21X1 _12738_ (
    .A(multiplier_0.reshi_5_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04864_)
  );
  NAND2X1 _12739_ (
    .A(_00121_),
    .B(_04839_),
    .Y(_04865_)
  );
  OAI21X1 _12740_ (
    .A(_04863_),
    .B(_04864_),
    .C(_04865_),
    .Y(_04417_)
  );
  XNOR2X1 _12741_ (
    .A(_04580_),
    .B(_04701_),
    .Y(_04866_)
  );
  OAI21X1 _12742_ (
    .A(multiplier_0.reshi_6_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04867_)
  );
  AOI21X1 _12743_ (
    .A(_05095_),
    .B(_04866_),
    .C(_04867_),
    .Y(_04868_)
  );
  AOI21X1 _12744_ (
    .A(_00122_),
    .B(_04839_),
    .C(_04868_),
    .Y(_04869_)
  );
  INVX1 _12745_ (
    .A(_04869_),
    .Y(_04418_)
  );
  XNOR2X1 _12746_ (
    .A(_04576_),
    .B(_04702_),
    .Y(_04870_)
  );
  AOI21X1 _12747_ (
    .A(_05095_),
    .B(_04870_),
    .C(_04843_),
    .Y(_04871_)
  );
  OAI21X1 _12748_ (
    .A(multiplier_0.reshi_7_ ),
    .B(_05095_),
    .C(_04871_),
    .Y(_04872_)
  );
  OAI21X1 _12749_ (
    .A(_05078_),
    .B(_04842_),
    .C(_04872_),
    .Y(_04419_)
  );
  XNOR2X1 _12750_ (
    .A(_04569_),
    .B(_04703_),
    .Y(_04873_)
  );
  AOI21X1 _12751_ (
    .A(_05095_),
    .B(_04873_),
    .C(_04843_),
    .Y(_04874_)
  );
  OAI21X1 _12752_ (
    .A(multiplier_0.reshi_8_ ),
    .B(_05095_),
    .C(_04874_),
    .Y(_04875_)
  );
  OAI21X1 _12753_ (
    .A(_04755_),
    .B(_04842_),
    .C(_04875_),
    .Y(_04420_)
  );
  NAND2X1 _12754_ (
    .A(_04561_),
    .B(_04562_),
    .Y(_04876_)
  );
  XNOR2X1 _12755_ (
    .A(_04704_),
    .B(_04876_),
    .Y(_04877_)
  );
  OAI21X1 _12756_ (
    .A(multiplier_0.reshi_9_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04878_)
  );
  INVX1 _12757_ (
    .A(_04878_),
    .Y(_04879_)
  );
  OAI21X1 _12758_ (
    .A(_05094_),
    .B(_04877_),
    .C(_04879_),
    .Y(_04880_)
  );
  OAI21X1 _12759_ (
    .A(_04757_),
    .B(_04842_),
    .C(_04880_),
    .Y(_04421_)
  );
  XOR2X1 _12760_ (
    .A(_04557_),
    .B(_04705_),
    .Y(_04881_)
  );
  OAI21X1 _12761_ (
    .A(multiplier_0.reshi_10_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04882_)
  );
  INVX1 _12762_ (
    .A(_04882_),
    .Y(_04883_)
  );
  OAI21X1 _12763_ (
    .A(_05094_),
    .B(_04881_),
    .C(_04883_),
    .Y(_04884_)
  );
  OAI21X1 _12764_ (
    .A(_04759_),
    .B(_04842_),
    .C(_04884_),
    .Y(_04407_)
  );
  NAND2X1 _12765_ (
    .A(_04550_),
    .B(_04551_),
    .Y(_04885_)
  );
  XOR2X1 _12766_ (
    .A(_04706_),
    .B(_04885_),
    .Y(_04886_)
  );
  AOI21X1 _12767_ (
    .A(_05095_),
    .B(_04886_),
    .C(_04843_),
    .Y(_04887_)
  );
  OAI21X1 _12768_ (
    .A(multiplier_0.reshi_11_ ),
    .B(_05095_),
    .C(_04887_),
    .Y(_04888_)
  );
  OAI21X1 _12769_ (
    .A(_04761_),
    .B(_04842_),
    .C(_04888_),
    .Y(_04408_)
  );
  XOR2X1 _12770_ (
    .A(_04546_),
    .B(_04707_),
    .Y(_04889_)
  );
  OAI21X1 _12771_ (
    .A(multiplier_0.reshi_12_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04890_)
  );
  INVX1 _12772_ (
    .A(_04890_),
    .Y(_04891_)
  );
  OAI21X1 _12773_ (
    .A(_05094_),
    .B(_04889_),
    .C(_04891_),
    .Y(_04892_)
  );
  OAI21X1 _12774_ (
    .A(_04763_),
    .B(_04842_),
    .C(_04892_),
    .Y(_04409_)
  );
  NAND2X1 _12775_ (
    .A(_04539_),
    .B(_04541_),
    .Y(_04893_)
  );
  XNOR2X1 _12776_ (
    .A(_04708_),
    .B(_04893_),
    .Y(_04894_)
  );
  OAI21X1 _12777_ (
    .A(multiplier_0.reshi_13_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04895_)
  );
  INVX1 _12778_ (
    .A(_04895_),
    .Y(_04896_)
  );
  OAI21X1 _12779_ (
    .A(_05094_),
    .B(_04894_),
    .C(_04896_),
    .Y(_04897_)
  );
  OAI21X1 _12780_ (
    .A(_04765_),
    .B(_04842_),
    .C(_04897_),
    .Y(_04410_)
  );
  XNOR2X1 _12781_ (
    .A(_04535_),
    .B(_04709_),
    .Y(_04898_)
  );
  OAI21X1 _12782_ (
    .A(multiplier_0.reshi_14_ ),
    .B(_05095_),
    .C(_04841_),
    .Y(_04899_)
  );
  AOI21X1 _12783_ (
    .A(_05095_),
    .B(_04898_),
    .C(_04899_),
    .Y(_04900_)
  );
  INVX1 _12784_ (
    .A(_04900_),
    .Y(_04901_)
  );
  OAI21X1 _12785_ (
    .A(_04767_),
    .B(_04842_),
    .C(_04901_),
    .Y(_04411_)
  );
  AOI21X1 _12786_ (
    .A(_05095_),
    .B(_04712_),
    .C(_04843_),
    .Y(_04902_)
  );
  OAI21X1 _12787_ (
    .A(multiplier_0.reshi_15_ ),
    .B(_05095_),
    .C(_04902_),
    .Y(_04903_)
  );
  OAI21X1 _12788_ (
    .A(_04769_),
    .B(_04842_),
    .C(_04903_),
    .Y(_04412_)
  );
  OR2X1 _12789_ (
    .A(_00102_),
    .B(_04723_),
    .Y(_04904_)
  );
  MUX2X1 _12790_ (
    .A(multiplier_0.acc_sel ),
    .B(_00101_),
    .S(_04904_),
    .Y(_04905_)
  );
  INVX1 _12791_ (
    .A(_04905_),
    .Y(_04373_)
  );
  MUX2X1 _12792_ (
    .A(multiplier_0.sign_sel ),
    .B(_00097_),
    .S(_04904_),
    .Y(_04906_)
  );
  INVX1 _12793_ (
    .A(_04906_),
    .Y(_04438_)
  );
  MUX2X1 _12794_ (
    .A(multiplier_0.op1_0_ ),
    .B(_00110_),
    .S(_04904_),
    .Y(_04907_)
  );
  INVX1 _12795_ (
    .A(_04907_),
    .Y(_04374_)
  );
  MUX2X1 _12796_ (
    .A(multiplier_0.op1_1_ ),
    .B(_00117_),
    .S(_04904_),
    .Y(_04908_)
  );
  INVX1 _12797_ (
    .A(_04908_),
    .Y(_04381_)
  );
  MUX2X1 _12798_ (
    .A(multiplier_0.op1_2_ ),
    .B(_00118_),
    .S(_04904_),
    .Y(_04909_)
  );
  INVX1 _12799_ (
    .A(_04909_),
    .Y(_04382_)
  );
  MUX2X1 _12800_ (
    .A(multiplier_0.op1_3_ ),
    .B(_00119_),
    .S(_04904_),
    .Y(_04910_)
  );
  INVX1 _12801_ (
    .A(_04910_),
    .Y(_04383_)
  );
  MUX2X1 _12802_ (
    .A(multiplier_0.op1_4_ ),
    .B(_00120_),
    .S(_04904_),
    .Y(_04911_)
  );
  INVX1 _12803_ (
    .A(_04911_),
    .Y(_04384_)
  );
  MUX2X1 _12804_ (
    .A(multiplier_0.op1_5_ ),
    .B(_00121_),
    .S(_04904_),
    .Y(_04912_)
  );
  INVX1 _12805_ (
    .A(_04912_),
    .Y(_04385_)
  );
  MUX2X1 _12806_ (
    .A(multiplier_0.op1_6_ ),
    .B(_00122_),
    .S(_04904_),
    .Y(_04913_)
  );
  INVX1 _12807_ (
    .A(_04913_),
    .Y(_04386_)
  );
  MUX2X1 _12808_ (
    .A(multiplier_0.op1_7_ ),
    .B(_00123_),
    .S(_04904_),
    .Y(_04914_)
  );
  INVX1 _12809_ (
    .A(_04914_),
    .Y(_04387_)
  );
  OAI21X1 _12810_ (
    .A(_00102_),
    .B(_05092_),
    .C(multiplier_0.op1_8_ ),
    .Y(_04915_)
  );
  OAI21X1 _12811_ (
    .A(_04755_),
    .B(_04904_),
    .C(_04915_),
    .Y(_04388_)
  );
  OAI21X1 _12812_ (
    .A(_00102_),
    .B(_05092_),
    .C(multiplier_0.op1_9_ ),
    .Y(_04916_)
  );
  OAI21X1 _12813_ (
    .A(_04757_),
    .B(_04904_),
    .C(_04916_),
    .Y(_04389_)
  );
  OAI21X1 _12814_ (
    .A(_00102_),
    .B(_05092_),
    .C(multiplier_0.op1_10_ ),
    .Y(_04917_)
  );
  OAI21X1 _12815_ (
    .A(_04759_),
    .B(_04904_),
    .C(_04917_),
    .Y(_04375_)
  );
  OAI21X1 _12816_ (
    .A(_00102_),
    .B(_05092_),
    .C(multiplier_0.op1_11_ ),
    .Y(_04918_)
  );
  OAI21X1 _12817_ (
    .A(_04761_),
    .B(_04904_),
    .C(_04918_),
    .Y(_04376_)
  );
  OAI21X1 _12818_ (
    .A(_00102_),
    .B(_05092_),
    .C(multiplier_0.op1_12_ ),
    .Y(_04919_)
  );
  OAI21X1 _12819_ (
    .A(_04763_),
    .B(_04904_),
    .C(_04919_),
    .Y(_04377_)
  );
  OAI21X1 _12820_ (
    .A(_00102_),
    .B(_05092_),
    .C(multiplier_0.op1_13_ ),
    .Y(_04920_)
  );
  OAI21X1 _12821_ (
    .A(_04765_),
    .B(_04904_),
    .C(_04920_),
    .Y(_04378_)
  );
  OAI21X1 _12822_ (
    .A(_00102_),
    .B(_05092_),
    .C(multiplier_0.op1_14_ ),
    .Y(_04921_)
  );
  OAI21X1 _12823_ (
    .A(_04767_),
    .B(_04904_),
    .C(_04921_),
    .Y(_04379_)
  );
  OAI21X1 _12824_ (
    .A(_00102_),
    .B(_05092_),
    .C(multiplier_0.op1_15_ ),
    .Y(_04922_)
  );
  OAI21X1 _12825_ (
    .A(_04769_),
    .B(_04904_),
    .C(_04922_),
    .Y(_04380_)
  );
  NOR3X1 _12826_ (
    .A(_05048_),
    .B(_04713_),
    .C(_04715_),
    .Y(_04923_)
  );
  NAND2X1 _12827_ (
    .A(_05090_),
    .B(_05091_),
    .Y(_04924_)
  );
  NAND3X1 _12828_ (
    .A(_00101_),
    .B(_05090_),
    .C(_05091_),
    .Y(_04925_)
  );
  NOR2X1 _12829_ (
    .A(_04772_),
    .B(_04925_),
    .Y(_04926_)
  );
  OAI21X1 _12830_ (
    .A(multiplier_0.sumext_0_ ),
    .B(multiplier_0.cycle_1_ ),
    .C(_04926_),
    .Y(_04927_)
  );
  NOR2X1 _12831_ (
    .A(_05079_),
    .B(_04925_),
    .Y(_04928_)
  );
  OAI21X1 _12832_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_0_ ),
    .C(_04928_),
    .Y(_04929_)
  );
  AOI21X1 _12833_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04837_),
    .C(_04929_),
    .Y(_04930_)
  );
  NOR2X1 _12834_ (
    .A(_04773_),
    .B(_04924_),
    .Y(_04931_)
  );
  OR2X1 _12835_ (
    .A(_04773_),
    .B(_04924_),
    .Y(_04932_)
  );
  NAND2X1 _12836_ (
    .A(_04771_),
    .B(_04931_),
    .Y(_04933_)
  );
  NOR2X1 _12837_ (
    .A(_05080_),
    .B(_04924_),
    .Y(_04934_)
  );
  NOR2X1 _12838_ (
    .A(_00102_),
    .B(_04924_),
    .Y(_04935_)
  );
  AOI22X1 _12839_ (
    .A(multiplier_0.op2_0_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_0_ ),
    .Y(_04936_)
  );
  NAND2X1 _12840_ (
    .A(_04933_),
    .B(_04936_),
    .Y(_04937_)
  );
  NOR2X1 _12841_ (
    .A(_04930_),
    .B(_04937_),
    .Y(_04938_)
  );
  OAI21X1 _12842_ (
    .A(_04923_),
    .B(_04927_),
    .C(_04938_),
    .Y(multiplier_0.per_dout_0_ )
  );
  OAI21X1 _12843_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.sumext_10_ ),
    .C(_04926_),
    .Y(_04939_)
  );
  INVX1 _12844_ (
    .A(_04939_),
    .Y(_04940_)
  );
  OAI21X1 _12845_ (
    .A(_05048_),
    .B(_04713_),
    .C(_04940_),
    .Y(_04941_)
  );
  OAI21X1 _12846_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_1_ ),
    .C(_04928_),
    .Y(_04942_)
  );
  AOI21X1 _12847_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04846_),
    .C(_04942_),
    .Y(_04943_)
  );
  NAND2X1 _12848_ (
    .A(_04783_),
    .B(_04931_),
    .Y(_04944_)
  );
  AOI22X1 _12849_ (
    .A(multiplier_0.op2_1_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_1_ ),
    .Y(_04945_)
  );
  NAND2X1 _12850_ (
    .A(_04944_),
    .B(_04945_),
    .Y(_04946_)
  );
  NOR2X1 _12851_ (
    .A(_04943_),
    .B(_04946_),
    .Y(_04947_)
  );
  NAND2X1 _12852_ (
    .A(_04941_),
    .B(_04947_),
    .Y(multiplier_0.per_dout_1_ )
  );
  OAI21X1 _12853_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_2_ ),
    .C(_04928_),
    .Y(_04948_)
  );
  AOI21X1 _12854_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04850_),
    .C(_04948_),
    .Y(_04949_)
  );
  NAND2X1 _12855_ (
    .A(_04787_),
    .B(_04931_),
    .Y(_04950_)
  );
  AOI22X1 _12856_ (
    .A(multiplier_0.op2_2_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_2_ ),
    .Y(_04951_)
  );
  NAND2X1 _12857_ (
    .A(_04950_),
    .B(_04951_),
    .Y(_04952_)
  );
  NOR2X1 _12858_ (
    .A(_04949_),
    .B(_04952_),
    .Y(_04953_)
  );
  NAND2X1 _12859_ (
    .A(_04941_),
    .B(_04953_),
    .Y(multiplier_0.per_dout_2_ )
  );
  OAI21X1 _12860_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_3_ ),
    .C(_04928_),
    .Y(_04954_)
  );
  AOI21X1 _12861_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04854_),
    .C(_04954_),
    .Y(_04955_)
  );
  NAND2X1 _12862_ (
    .A(_04791_),
    .B(_04931_),
    .Y(_04956_)
  );
  AOI22X1 _12863_ (
    .A(multiplier_0.op2_3_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_3_ ),
    .Y(_04957_)
  );
  NAND2X1 _12864_ (
    .A(_04956_),
    .B(_04957_),
    .Y(_04958_)
  );
  NOR2X1 _12865_ (
    .A(_04955_),
    .B(_04958_),
    .Y(_04959_)
  );
  NAND2X1 _12866_ (
    .A(_04941_),
    .B(_04959_),
    .Y(multiplier_0.per_dout_3_ )
  );
  OAI21X1 _12867_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_4_ ),
    .C(_04928_),
    .Y(_04960_)
  );
  AOI21X1 _12868_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04858_),
    .C(_04960_),
    .Y(_04961_)
  );
  AOI22X1 _12869_ (
    .A(multiplier_0.op2_4_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_4_ ),
    .Y(_04962_)
  );
  OAI21X1 _12870_ (
    .A(_04795_),
    .B(_04932_),
    .C(_04962_),
    .Y(_04963_)
  );
  NOR2X1 _12871_ (
    .A(_04961_),
    .B(_04963_),
    .Y(_04964_)
  );
  NAND2X1 _12872_ (
    .A(_04941_),
    .B(_04964_),
    .Y(multiplier_0.per_dout_4_ )
  );
  NOR2X1 _12873_ (
    .A(_05048_),
    .B(_04862_),
    .Y(_04965_)
  );
  OAI21X1 _12874_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_5_ ),
    .C(_04928_),
    .Y(_04966_)
  );
  NOR2X1 _12875_ (
    .A(_04965_),
    .B(_04966_),
    .Y(_04967_)
  );
  AOI22X1 _12876_ (
    .A(multiplier_0.op2_5_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_5_ ),
    .Y(_04968_)
  );
  OAI21X1 _12877_ (
    .A(_04799_),
    .B(_04932_),
    .C(_04968_),
    .Y(_04969_)
  );
  NOR2X1 _12878_ (
    .A(_04967_),
    .B(_04969_),
    .Y(_04970_)
  );
  NAND2X1 _12879_ (
    .A(_04941_),
    .B(_04970_),
    .Y(multiplier_0.per_dout_5_ )
  );
  OAI21X1 _12880_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_6_ ),
    .C(_04928_),
    .Y(_04971_)
  );
  AOI21X1 _12881_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04866_),
    .C(_04971_),
    .Y(_04972_)
  );
  NAND2X1 _12882_ (
    .A(_04803_),
    .B(_04931_),
    .Y(_04973_)
  );
  AOI22X1 _12883_ (
    .A(multiplier_0.op2_6_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_6_ ),
    .Y(_04974_)
  );
  NAND2X1 _12884_ (
    .A(_04973_),
    .B(_04974_),
    .Y(_04975_)
  );
  NOR2X1 _12885_ (
    .A(_04972_),
    .B(_04975_),
    .Y(_04976_)
  );
  NAND2X1 _12886_ (
    .A(_04941_),
    .B(_04976_),
    .Y(multiplier_0.per_dout_6_ )
  );
  OAI21X1 _12887_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_7_ ),
    .C(_04928_),
    .Y(_04977_)
  );
  AOI21X1 _12888_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04870_),
    .C(_04977_),
    .Y(_04978_)
  );
  AOI22X1 _12889_ (
    .A(multiplier_0.op2_7_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_7_ ),
    .Y(_04979_)
  );
  OAI21X1 _12890_ (
    .A(_04807_),
    .B(_04932_),
    .C(_04979_),
    .Y(_04980_)
  );
  NOR2X1 _12891_ (
    .A(_04978_),
    .B(_04980_),
    .Y(_04981_)
  );
  NAND2X1 _12892_ (
    .A(_04941_),
    .B(_04981_),
    .Y(multiplier_0.per_dout_7_ )
  );
  OAI21X1 _12893_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_8_ ),
    .C(_04928_),
    .Y(_04982_)
  );
  AOI21X1 _12894_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04873_),
    .C(_04982_),
    .Y(_04983_)
  );
  AND2X1 _12895_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04809_),
    .Y(_04984_)
  );
  OAI21X1 _12896_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_8_ ),
    .C(_04931_),
    .Y(_04985_)
  );
  AOI22X1 _12897_ (
    .A(multiplier_0.op2_8_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_8_ ),
    .Y(_04986_)
  );
  OAI21X1 _12898_ (
    .A(_04984_),
    .B(_04985_),
    .C(_04986_),
    .Y(_04987_)
  );
  NOR2X1 _12899_ (
    .A(_04983_),
    .B(_04987_),
    .Y(_04988_)
  );
  NAND2X1 _12900_ (
    .A(_04941_),
    .B(_04988_),
    .Y(multiplier_0.per_dout_8_ )
  );
  NOR2X1 _12901_ (
    .A(_05048_),
    .B(_04877_),
    .Y(_04989_)
  );
  OAI21X1 _12902_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_9_ ),
    .C(_04928_),
    .Y(_04990_)
  );
  NOR2X1 _12903_ (
    .A(_04989_),
    .B(_04990_),
    .Y(_04991_)
  );
  AND2X1 _12904_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04812_),
    .Y(_04992_)
  );
  OAI21X1 _12905_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_9_ ),
    .C(_04931_),
    .Y(_04993_)
  );
  AOI22X1 _12906_ (
    .A(multiplier_0.op2_9_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_9_ ),
    .Y(_04994_)
  );
  OAI21X1 _12907_ (
    .A(_04992_),
    .B(_04993_),
    .C(_04994_),
    .Y(_04995_)
  );
  NOR2X1 _12908_ (
    .A(_04991_),
    .B(_04995_),
    .Y(_04996_)
  );
  NAND2X1 _12909_ (
    .A(_04941_),
    .B(_04996_),
    .Y(multiplier_0.per_dout_9_ )
  );
  NOR2X1 _12910_ (
    .A(_05048_),
    .B(_04881_),
    .Y(_04997_)
  );
  OAI21X1 _12911_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_10_ ),
    .C(_04928_),
    .Y(_04998_)
  );
  NOR2X1 _12912_ (
    .A(_04997_),
    .B(_04998_),
    .Y(_04999_)
  );
  AND2X1 _12913_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04816_),
    .Y(_05000_)
  );
  OAI21X1 _12914_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_10_ ),
    .C(_04931_),
    .Y(_05001_)
  );
  AOI22X1 _12915_ (
    .A(multiplier_0.op2_10_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_10_ ),
    .Y(_05002_)
  );
  OAI21X1 _12916_ (
    .A(_05000_),
    .B(_05001_),
    .C(_05002_),
    .Y(_05003_)
  );
  NOR2X1 _12917_ (
    .A(_04999_),
    .B(_05003_),
    .Y(_05004_)
  );
  NAND2X1 _12918_ (
    .A(_04941_),
    .B(_05004_),
    .Y(multiplier_0.per_dout_10_ )
  );
  OAI21X1 _12919_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_11_ ),
    .C(_04928_),
    .Y(_05005_)
  );
  AOI21X1 _12920_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04886_),
    .C(_05005_),
    .Y(_05006_)
  );
  AND2X1 _12921_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04819_),
    .Y(_05007_)
  );
  OAI21X1 _12922_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_11_ ),
    .C(_04931_),
    .Y(_05008_)
  );
  AOI22X1 _12923_ (
    .A(multiplier_0.op2_11_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_11_ ),
    .Y(_05009_)
  );
  OAI21X1 _12924_ (
    .A(_05007_),
    .B(_05008_),
    .C(_05009_),
    .Y(_05010_)
  );
  NOR2X1 _12925_ (
    .A(_05006_),
    .B(_05010_),
    .Y(_05011_)
  );
  NAND2X1 _12926_ (
    .A(_04941_),
    .B(_05011_),
    .Y(multiplier_0.per_dout_11_ )
  );
  NOR2X1 _12927_ (
    .A(_05048_),
    .B(_04889_),
    .Y(_05012_)
  );
  OAI21X1 _12928_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_12_ ),
    .C(_04928_),
    .Y(_05013_)
  );
  NOR2X1 _12929_ (
    .A(_05012_),
    .B(_05013_),
    .Y(_05014_)
  );
  AND2X1 _12930_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04822_),
    .Y(_05015_)
  );
  OAI21X1 _12931_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_12_ ),
    .C(_04931_),
    .Y(_05016_)
  );
  AOI22X1 _12932_ (
    .A(multiplier_0.op2_12_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_12_ ),
    .Y(_05017_)
  );
  OAI21X1 _12933_ (
    .A(_05015_),
    .B(_05016_),
    .C(_05017_),
    .Y(_05018_)
  );
  NOR2X1 _12934_ (
    .A(_05014_),
    .B(_05018_),
    .Y(_05019_)
  );
  NAND2X1 _12935_ (
    .A(_04941_),
    .B(_05019_),
    .Y(multiplier_0.per_dout_12_ )
  );
  NOR2X1 _12936_ (
    .A(_05048_),
    .B(_04894_),
    .Y(_05020_)
  );
  OAI21X1 _12937_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_13_ ),
    .C(_04928_),
    .Y(_05021_)
  );
  NOR2X1 _12938_ (
    .A(_05020_),
    .B(_05021_),
    .Y(_05022_)
  );
  AND2X1 _12939_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04826_),
    .Y(_05023_)
  );
  OAI21X1 _12940_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_13_ ),
    .C(_04931_),
    .Y(_05024_)
  );
  AOI22X1 _12941_ (
    .A(multiplier_0.op2_13_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_13_ ),
    .Y(_05025_)
  );
  OAI21X1 _12942_ (
    .A(_05023_),
    .B(_05024_),
    .C(_05025_),
    .Y(_05026_)
  );
  NOR2X1 _12943_ (
    .A(_05022_),
    .B(_05026_),
    .Y(_05027_)
  );
  NAND2X1 _12944_ (
    .A(_04941_),
    .B(_05027_),
    .Y(multiplier_0.per_dout_13_ )
  );
  OAI21X1 _12945_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_14_ ),
    .C(_04928_),
    .Y(_05028_)
  );
  AOI21X1 _12946_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04898_),
    .C(_05028_),
    .Y(_05029_)
  );
  AND2X1 _12947_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04830_),
    .Y(_05030_)
  );
  OAI21X1 _12948_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_14_ ),
    .C(_04931_),
    .Y(_05031_)
  );
  AOI22X1 _12949_ (
    .A(multiplier_0.op2_14_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_14_ ),
    .Y(_05032_)
  );
  OAI21X1 _12950_ (
    .A(_05030_),
    .B(_05031_),
    .C(_05032_),
    .Y(_05033_)
  );
  NOR2X1 _12951_ (
    .A(_05029_),
    .B(_05033_),
    .Y(_05034_)
  );
  NAND2X1 _12952_ (
    .A(_04941_),
    .B(_05034_),
    .Y(multiplier_0.per_dout_14_ )
  );
  OAI21X1 _12953_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reshi_15_ ),
    .C(_04928_),
    .Y(_05035_)
  );
  AOI21X1 _12954_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04712_),
    .C(_05035_),
    .Y(_05036_)
  );
  AND2X1 _12955_ (
    .A(multiplier_0.cycle_1_ ),
    .B(_04833_),
    .Y(_05037_)
  );
  OAI21X1 _12956_ (
    .A(multiplier_0.cycle_1_ ),
    .B(multiplier_0.reslo_15_ ),
    .C(_04931_),
    .Y(_05038_)
  );
  AOI22X1 _12957_ (
    .A(multiplier_0.op2_15_ ),
    .B(_04934_),
    .C(_04935_),
    .D(multiplier_0.op1_15_ ),
    .Y(_05039_)
  );
  OAI21X1 _12958_ (
    .A(_05037_),
    .B(_05038_),
    .C(_05039_),
    .Y(_05040_)
  );
  NOR2X1 _12959_ (
    .A(_05036_),
    .B(_05040_),
    .Y(_05041_)
  );
  NAND2X1 _12960_ (
    .A(_04941_),
    .B(_05041_),
    .Y(multiplier_0.per_dout_15_ )
  );
  DFFSR _12961_ (
    .CLK(dco_clk),
    .D(multiplier_0.op2_wr ),
    .Q(multiplier_0.cycle_0_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12962_ (
    .CLK(dco_clk),
    .D(multiplier_0.cycle_0_ ),
    .Q(multiplier_0.cycle_1_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12963_ (
    .CLK(dco_clk),
    .D(_04373_),
    .Q(multiplier_0.acc_sel ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12964_ (
    .CLK(dco_clk),
    .D(_04438_),
    .Q(multiplier_0.sign_sel ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12965_ (
    .CLK(dco_clk),
    .D(_04439_),
    .Q(multiplier_0.sumext_0_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12966_ (
    .CLK(dco_clk),
    .D(_04440_),
    .Q(multiplier_0.sumext_10_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12967_ (
    .CLK(dco_clk),
    .D(_04406_),
    .Q(multiplier_0.reshi_0_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12968_ (
    .CLK(dco_clk),
    .D(_04413_),
    .Q(multiplier_0.reshi_1_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12969_ (
    .CLK(dco_clk),
    .D(_04414_),
    .Q(multiplier_0.reshi_2_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12970_ (
    .CLK(dco_clk),
    .D(_04415_),
    .Q(multiplier_0.reshi_3_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12971_ (
    .CLK(dco_clk),
    .D(_04416_),
    .Q(multiplier_0.reshi_4_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12972_ (
    .CLK(dco_clk),
    .D(_04417_),
    .Q(multiplier_0.reshi_5_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12973_ (
    .CLK(dco_clk),
    .D(_04418_),
    .Q(multiplier_0.reshi_6_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12974_ (
    .CLK(dco_clk),
    .D(_04419_),
    .Q(multiplier_0.reshi_7_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12975_ (
    .CLK(dco_clk),
    .D(_04420_),
    .Q(multiplier_0.reshi_8_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12976_ (
    .CLK(dco_clk),
    .D(_04421_),
    .Q(multiplier_0.reshi_9_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12977_ (
    .CLK(dco_clk),
    .D(_04407_),
    .Q(multiplier_0.reshi_10_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12978_ (
    .CLK(dco_clk),
    .D(_04408_),
    .Q(multiplier_0.reshi_11_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12979_ (
    .CLK(dco_clk),
    .D(_04409_),
    .Q(multiplier_0.reshi_12_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12980_ (
    .CLK(dco_clk),
    .D(_04410_),
    .Q(multiplier_0.reshi_13_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12981_ (
    .CLK(dco_clk),
    .D(_04411_),
    .Q(multiplier_0.reshi_14_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12982_ (
    .CLK(dco_clk),
    .D(_04412_),
    .Q(multiplier_0.reshi_15_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12983_ (
    .CLK(dco_clk),
    .D(_04422_),
    .Q(multiplier_0.reslo_0_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12984_ (
    .CLK(dco_clk),
    .D(_04429_),
    .Q(multiplier_0.reslo_1_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12985_ (
    .CLK(dco_clk),
    .D(_04430_),
    .Q(multiplier_0.reslo_2_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12986_ (
    .CLK(dco_clk),
    .D(_04431_),
    .Q(multiplier_0.reslo_3_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12987_ (
    .CLK(dco_clk),
    .D(_04432_),
    .Q(multiplier_0.reslo_4_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12988_ (
    .CLK(dco_clk),
    .D(_04433_),
    .Q(multiplier_0.reslo_5_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12989_ (
    .CLK(dco_clk),
    .D(_04434_),
    .Q(multiplier_0.reslo_6_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12990_ (
    .CLK(dco_clk),
    .D(_04435_),
    .Q(multiplier_0.reslo_7_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12991_ (
    .CLK(dco_clk),
    .D(_04436_),
    .Q(multiplier_0.reslo_8_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12992_ (
    .CLK(dco_clk),
    .D(_04437_),
    .Q(multiplier_0.reslo_9_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12993_ (
    .CLK(dco_clk),
    .D(_04423_),
    .Q(multiplier_0.reslo_10_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12994_ (
    .CLK(dco_clk),
    .D(_04424_),
    .Q(multiplier_0.reslo_11_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12995_ (
    .CLK(dco_clk),
    .D(_04425_),
    .Q(multiplier_0.reslo_12_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12996_ (
    .CLK(dco_clk),
    .D(_04426_),
    .Q(multiplier_0.reslo_13_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12997_ (
    .CLK(dco_clk),
    .D(_04427_),
    .Q(multiplier_0.reslo_14_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12998_ (
    .CLK(dco_clk),
    .D(_04428_),
    .Q(multiplier_0.reslo_15_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _12999_ (
    .CLK(dco_clk),
    .D(_04390_),
    .Q(multiplier_0.op2_0_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13000_ (
    .CLK(dco_clk),
    .D(_04397_),
    .Q(multiplier_0.op2_1_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13001_ (
    .CLK(dco_clk),
    .D(_04398_),
    .Q(multiplier_0.op2_2_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13002_ (
    .CLK(dco_clk),
    .D(_04399_),
    .Q(multiplier_0.op2_3_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13003_ (
    .CLK(dco_clk),
    .D(_04400_),
    .Q(multiplier_0.op2_4_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13004_ (
    .CLK(dco_clk),
    .D(_04401_),
    .Q(multiplier_0.op2_5_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13005_ (
    .CLK(dco_clk),
    .D(_04402_),
    .Q(multiplier_0.op2_6_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13006_ (
    .CLK(dco_clk),
    .D(_04403_),
    .Q(multiplier_0.op2_7_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13007_ (
    .CLK(dco_clk),
    .D(_04404_),
    .Q(multiplier_0.op2_8_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13008_ (
    .CLK(dco_clk),
    .D(_04405_),
    .Q(multiplier_0.op2_9_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13009_ (
    .CLK(dco_clk),
    .D(_04391_),
    .Q(multiplier_0.op2_10_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13010_ (
    .CLK(dco_clk),
    .D(_04392_),
    .Q(multiplier_0.op2_11_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13011_ (
    .CLK(dco_clk),
    .D(_04393_),
    .Q(multiplier_0.op2_12_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13012_ (
    .CLK(dco_clk),
    .D(_04394_),
    .Q(multiplier_0.op2_13_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13013_ (
    .CLK(dco_clk),
    .D(_04395_),
    .Q(multiplier_0.op2_14_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13014_ (
    .CLK(dco_clk),
    .D(_04396_),
    .Q(multiplier_0.op2_15_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13015_ (
    .CLK(dco_clk),
    .D(_04374_),
    .Q(multiplier_0.op1_0_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13016_ (
    .CLK(dco_clk),
    .D(_04381_),
    .Q(multiplier_0.op1_1_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13017_ (
    .CLK(dco_clk),
    .D(_04382_),
    .Q(multiplier_0.op1_2_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13018_ (
    .CLK(dco_clk),
    .D(_04383_),
    .Q(multiplier_0.op1_3_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13019_ (
    .CLK(dco_clk),
    .D(_04384_),
    .Q(multiplier_0.op1_4_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13020_ (
    .CLK(dco_clk),
    .D(_04385_),
    .Q(multiplier_0.op1_5_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13021_ (
    .CLK(dco_clk),
    .D(_04386_),
    .Q(multiplier_0.op1_6_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13022_ (
    .CLK(dco_clk),
    .D(_04387_),
    .Q(multiplier_0.op1_7_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13023_ (
    .CLK(dco_clk),
    .D(_04388_),
    .Q(multiplier_0.op1_8_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13024_ (
    .CLK(dco_clk),
    .D(_04389_),
    .Q(multiplier_0.op1_9_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13025_ (
    .CLK(dco_clk),
    .D(_04375_),
    .Q(multiplier_0.op1_10_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13026_ (
    .CLK(dco_clk),
    .D(_04376_),
    .Q(multiplier_0.op1_11_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13027_ (
    .CLK(dco_clk),
    .D(_04377_),
    .Q(multiplier_0.op1_12_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13028_ (
    .CLK(dco_clk),
    .D(_04378_),
    .Q(multiplier_0.op1_13_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13029_ (
    .CLK(dco_clk),
    .D(_04379_),
    .Q(multiplier_0.op1_14_ ),
    .R(_04441_),
    .S(1'h1)
  );
  DFFSR _13030_ (
    .CLK(dco_clk),
    .D(_04380_),
    .Q(multiplier_0.op1_15_ ),
    .R(_04441_),
    .S(1'h1)
  );
  INVX1 _13031_ (
    .A(_00097_),
    .Y(_05857_)
  );
  INVX1 _13032_ (
    .A(_00101_),
    .Y(_05858_)
  );
  INVX1 _13033_ (
    .A(_00100_),
    .Y(_05859_)
  );
  INVX1 _13034_ (
    .A(_00126_),
    .Y(_05860_)
  );
  INVX1 _13035_ (
    .A(_00110_),
    .Y(_05861_)
  );
  INVX1 _13036_ (
    .A(sfr_0.ie1_0_ ),
    .Y(_05862_)
  );
  INVX1 _13037_ (
    .A(1'h0),
    .Y(_05863_)
  );
  INVX1 _13038_ (
    .A(1'h0),
    .Y(_05864_)
  );
  INVX1 _13039_ (
    .A(1'h0),
    .Y(_05865_)
  );
  INVX1 _13040_ (
    .A(1'h0),
    .Y(_05866_)
  );
  INVX1 _13041_ (
    .A(sfr_0.ifg1_0_ ),
    .Y(_05867_)
  );
  INVX1 _13042_ (
    .A(_00162_),
    .Y(_05850_)
  );
  NOR2X1 _13043_ (
    .A(_00097_),
    .B(_00101_),
    .Y(_05868_)
  );
  INVX1 _13044_ (
    .A(_05868_),
    .Y(_05869_)
  );
  NOR2X1 _13045_ (
    .A(_00102_),
    .B(_05869_),
    .Y(_05870_)
  );
  NOR2X1 _13046_ (
    .A(_00099_),
    .B(1'h0),
    .Y(_05871_)
  );
  OR2X1 _13047_ (
    .A(_00099_),
    .B(1'h0),
    .Y(_05872_)
  );
  NOR3X1 _13048_ (
    .A(_00100_),
    .B(_05860_),
    .C(_05872_),
    .Y(_05873_)
  );
  NAND3X1 _13049_ (
    .A(_05859_),
    .B(_00126_),
    .C(_05871_),
    .Y(_05874_)
  );
  NOR2X1 _13050_ (
    .A(_00108_),
    .B(_00107_),
    .Y(_05875_)
  );
  NOR2X1 _13051_ (
    .A(_00098_),
    .B(_00109_),
    .Y(_05876_)
  );
  AND2X1 _13052_ (
    .A(_05875_),
    .B(_05876_),
    .Y(_05877_)
  );
  NAND2X1 _13053_ (
    .A(_05875_),
    .B(_05876_),
    .Y(_05878_)
  );
  NOR2X1 _13054_ (
    .A(_00104_),
    .B(_00103_),
    .Y(_05879_)
  );
  NOR2X1 _13055_ (
    .A(_00106_),
    .B(_00105_),
    .Y(_05880_)
  );
  AND2X1 _13056_ (
    .A(_05879_),
    .B(_05880_),
    .Y(_05881_)
  );
  NAND2X1 _13057_ (
    .A(_05879_),
    .B(_05880_),
    .Y(_05882_)
  );
  NOR3X1 _13058_ (
    .A(_05874_),
    .B(_05878_),
    .C(_05882_),
    .Y(_05883_)
  );
  NAND3X1 _13059_ (
    .A(_05873_),
    .B(_05877_),
    .C(_05881_),
    .Y(_05884_)
  );
  NAND3X1 _13060_ (
    .A(_00127_),
    .B(_05870_),
    .C(_05883_),
    .Y(_05885_)
  );
  MUX2X1 _13061_ (
    .A(_05862_),
    .B(_05861_),
    .S(_05885_),
    .Y(_05849_)
  );
  NOR2X1 _13062_ (
    .A(_05858_),
    .B(_00102_),
    .Y(_05886_)
  );
  NOR2X1 _13063_ (
    .A(_00127_),
    .B(_00128_),
    .Y(_05887_)
  );
  INVX1 _13064_ (
    .A(_05887_),
    .Y(_05888_)
  );
  NAND2X1 _13065_ (
    .A(_05883_),
    .B(_05887_),
    .Y(_05889_)
  );
  NAND3X1 _13066_ (
    .A(_05883_),
    .B(_05886_),
    .C(_05887_),
    .Y(_05890_)
  );
  AND2X1 _13067_ (
    .A(_00102_),
    .B(_05868_),
    .Y(_05891_)
  );
  NAND2X1 _13068_ (
    .A(_00102_),
    .B(_05868_),
    .Y(_05892_)
  );
  NOR3X1 _13069_ (
    .A(_05884_),
    .B(_05888_),
    .C(_05892_),
    .Y(_05893_)
  );
  NAND3X1 _13070_ (
    .A(_05883_),
    .B(_05887_),
    .C(_05891_),
    .Y(_05894_)
  );
  OAI22X1 _13071_ (
    .A(_00097_),
    .B(_05890_),
    .C(_05894_),
    .D(_05863_),
    .Y(per_dout_sfr_14_)
  );
  OAI22X1 _13072_ (
    .A(_05857_),
    .B(_05890_),
    .C(_05894_),
    .D(_05864_),
    .Y(per_dout_sfr_8_)
  );
  OAI22X1 _13073_ (
    .A(_05857_),
    .B(_05890_),
    .C(_05894_),
    .D(_05865_),
    .Y(per_dout_sfr_15_)
  );
  OAI22X1 _13074_ (
    .A(_00097_),
    .B(_05890_),
    .C(_05894_),
    .D(_05866_),
    .Y(per_dout_sfr_1_)
  );
  NAND2X1 _13075_ (
    .A(1'h0),
    .B(_05891_),
    .Y(_05851_)
  );
  OR2X1 _13076_ (
    .A(_05857_),
    .B(_00102_),
    .Y(_05852_)
  );
  OAI22X1 _13077_ (
    .A(_05858_),
    .B(_00102_),
    .C(_05867_),
    .D(_05852_),
    .Y(_05853_)
  );
  NOR2X1 _13078_ (
    .A(_00101_),
    .B(_05852_),
    .Y(_05854_)
  );
  AOI21X1 _13079_ (
    .A(sfr_0.ie1_0_ ),
    .B(_05870_),
    .C(_05853_),
    .Y(_05855_)
  );
  AOI21X1 _13080_ (
    .A(_05851_),
    .B(_05855_),
    .C(_05889_),
    .Y(per_dout_sfr_0_)
  );
  NAND3X1 _13081_ (
    .A(_00127_),
    .B(_05883_),
    .C(_05854_),
    .Y(_05856_)
  );
  NOR2X1 _13082_ (
    .A(_00110_),
    .B(_05856_),
    .Y(sfr_0.wdtifg_sw_clr )
  );
  NOR2X1 _13083_ (
    .A(_05861_),
    .B(_05856_),
    .Y(sfr_0.wdtifg_sw_set )
  );
  AND2X1 _13084_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_2_)
  );
  AND2X1 _13085_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_3_)
  );
  AND2X1 _13086_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_4_)
  );
  AND2X1 _13087_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_5_)
  );
  AND2X1 _13088_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_6_)
  );
  AND2X1 _13089_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_7_)
  );
  AND2X1 _13090_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_9_)
  );
  AND2X1 _13091_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_10_)
  );
  AND2X1 _13092_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_11_)
  );
  AND2X1 _13093_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_12_)
  );
  AND2X1 _13094_ (
    .A(1'h0),
    .B(_05893_),
    .Y(per_dout_sfr_13_)
  );
  DFFSR _13095_ (
    .CLK(dco_clk),
    .D(_05849_),
    .Q(sfr_0.ie1_0_ ),
    .R(_05850_),
    .S(1'h1)
  );
  INVX1 _13096_ (
    .A(_00048_),
    .Y(_05923_)
  );
  INVX1 _13097_ (
    .A(_00104_),
    .Y(_05924_)
  );
  INVX1 _13098_ (
    .A(_00106_),
    .Y(_05925_)
  );
  INVX1 _13099_ (
    .A(_00108_),
    .Y(_05926_)
  );
  INVX1 _13100_ (
    .A(1'h0),
    .Y(_05927_)
  );
  INVX1 _13101_ (
    .A(_00097_),
    .Y(_05928_)
  );
  INVX1 _13102_ (
    .A(watchdog_0.wdtcnt_6_ ),
    .Y(_05929_)
  );
  INVX1 _13103_ (
    .A(watchdog_0.wdtcnt_1_ ),
    .Y(_05930_)
  );
  INVX1 _13104_ (
    .A(watchdog_0.wdtctl_0_ ),
    .Y(_05931_)
  );
  INVX1 _13105_ (
    .A(watchdog_0.wdtctl_1_ ),
    .Y(_05932_)
  );
  INVX1 _13106_ (
    .A(watchdog_0.wdtcnt_9_ ),
    .Y(_05933_)
  );
  INVX1 _13107_ (
    .A(watchdog_0.wdtcnt_10_ ),
    .Y(_05934_)
  );
  INVX1 _13108_ (
    .A(_00119_),
    .Y(_05935_)
  );
  INVX1 _13109_ (
    .A(sfr_0.wdtifg_sw_clr ),
    .Y(_05936_)
  );
  INVX1 _13110_ (
    .A(sfr_0.wdtifg_sw_set ),
    .Y(_05937_)
  );
  INVX1 _13111_ (
    .A(clock_module_0.por ),
    .Y(_05921_)
  );
  INVX1 _13112_ (
    .A(_00162_),
    .Y(_05922_)
  );
  NAND2X1 _13113_ (
    .A(watchdog_0.wdtcnt_11_ ),
    .B(watchdog_0.wdtcnt_10_ ),
    .Y(_05938_)
  );
  NAND3X1 _13114_ (
    .A(watchdog_0.wdtcnt_12_ ),
    .B(watchdog_0.wdtcnt_11_ ),
    .C(watchdog_0.wdtcnt_10_ ),
    .Y(_05939_)
  );
  AND2X1 _13115_ (
    .A(watchdog_0.wdtcnt_3_ ),
    .B(watchdog_0.wdtcnt_2_ ),
    .Y(_05940_)
  );
  NAND2X1 _13116_ (
    .A(watchdog_0.wdtcnt_3_ ),
    .B(watchdog_0.wdtcnt_2_ ),
    .Y(_05941_)
  );
  AND2X1 _13117_ (
    .A(watchdog_0.wdtcnt_0_ ),
    .B(watchdog_0.wdtcnt_5_ ),
    .Y(_05942_)
  );
  NAND2X1 _13118_ (
    .A(watchdog_0.wdtcnt_0_ ),
    .B(watchdog_0.wdtcnt_5_ ),
    .Y(_05943_)
  );
  AND2X1 _13119_ (
    .A(watchdog_0.wdtcnt_4_ ),
    .B(watchdog_0.wdtcnt_1_ ),
    .Y(_05944_)
  );
  NAND2X1 _13120_ (
    .A(watchdog_0.wdtcnt_4_ ),
    .B(watchdog_0.wdtcnt_1_ ),
    .Y(_05945_)
  );
  NOR3X1 _13121_ (
    .A(_05941_),
    .B(_05943_),
    .C(_05945_),
    .Y(_05946_)
  );
  NAND3X1 _13122_ (
    .A(_05940_),
    .B(_05942_),
    .C(_05944_),
    .Y(_05947_)
  );
  NOR2X1 _13123_ (
    .A(_05929_),
    .B(_05947_),
    .Y(_05948_)
  );
  AND2X1 _13124_ (
    .A(watchdog_0.wdtcnt_7_ ),
    .B(watchdog_0.wdtcnt_8_ ),
    .Y(_05949_)
  );
  NAND2X1 _13125_ (
    .A(watchdog_0.wdtcnt_7_ ),
    .B(watchdog_0.wdtcnt_8_ ),
    .Y(_05950_)
  );
  NOR3X1 _13126_ (
    .A(_05929_),
    .B(_05947_),
    .C(_05950_),
    .Y(_05951_)
  );
  NAND3X1 _13127_ (
    .A(watchdog_0.wdtcnt_6_ ),
    .B(_05946_),
    .C(_05949_),
    .Y(_05952_)
  );
  NOR3X1 _13128_ (
    .A(_05933_),
    .B(_05939_),
    .C(_05952_),
    .Y(_05953_)
  );
  NAND3X1 _13129_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(watchdog_0.wdtcnt_14_ ),
    .C(_05953_),
    .Y(_05954_)
  );
  XOR2X1 _13130_ (
    .A(watchdog_0.wdtcnt_15_ ),
    .B(_05954_),
    .Y(_05955_)
  );
  XNOR2X1 _13131_ (
    .A(watchdog_0.wdtcnt_15_ ),
    .B(_05954_),
    .Y(_05956_)
  );
  NOR2X1 _13132_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(watchdog_0.wdtctl_1_ ),
    .Y(_05957_)
  );
  NAND2X1 _13133_ (
    .A(_05931_),
    .B(_05932_),
    .Y(_05958_)
  );
  XOR2X1 _13134_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(_05953_),
    .Y(_05959_)
  );
  XNOR2X1 _13135_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(_05953_),
    .Y(_05960_)
  );
  NAND2X1 _13136_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(watchdog_0.wdtctl_1_ ),
    .Y(_05961_)
  );
  NOR2X1 _13137_ (
    .A(watchdog_0.wdtcnt_9_ ),
    .B(_05951_),
    .Y(_05962_)
  );
  NAND2X1 _13138_ (
    .A(_05933_),
    .B(_05952_),
    .Y(_05963_)
  );
  AOI21X1 _13139_ (
    .A(watchdog_0.wdtcnt_9_ ),
    .B(_05951_),
    .C(_05932_),
    .Y(_05964_)
  );
  OAI21X1 _13140_ (
    .A(_05933_),
    .B(_05952_),
    .C(watchdog_0.wdtctl_1_ ),
    .Y(_05965_)
  );
  AOI22X1 _13141_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(watchdog_0.wdtctl_1_ ),
    .C(_05963_),
    .D(_05964_),
    .Y(_05966_)
  );
  OAI21X1 _13142_ (
    .A(_05962_),
    .B(_05965_),
    .C(_05961_),
    .Y(_05967_)
  );
  AOI21X1 _13143_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(_05959_),
    .C(_05967_),
    .Y(_05968_)
  );
  OAI21X1 _13144_ (
    .A(_05931_),
    .B(_05960_),
    .C(_05966_),
    .Y(_05969_)
  );
  AOI21X1 _13145_ (
    .A(_05956_),
    .B(_05957_),
    .C(_05969_),
    .Y(_05970_)
  );
  OAI21X1 _13146_ (
    .A(_05955_),
    .B(_05958_),
    .C(_05968_),
    .Y(_05971_)
  );
  OR2X1 _13147_ (
    .A(watchdog_0.wdtctl_7_ ),
    .B(_00049_),
    .Y(_05972_)
  );
  OR2X1 _13148_ (
    .A(_00163_),
    .B(watchdog_0.wdtctl_2_ ),
    .Y(_05973_)
  );
  AOI21X1 _13149_ (
    .A(_05923_),
    .B(watchdog_0.wdtctl_2_ ),
    .C(_05972_),
    .Y(_05974_)
  );
  AND2X1 _13150_ (
    .A(_05973_),
    .B(_05974_),
    .Y(_05975_)
  );
  OAI21X1 _13151_ (
    .A(_00163_),
    .B(watchdog_0.wdtctl_2_ ),
    .C(_05974_),
    .Y(_05976_)
  );
  OAI21X1 _13152_ (
    .A(watchdog_0.wdtcnt_6_ ),
    .B(_05946_),
    .C(_05975_),
    .Y(_05977_)
  );
  NOR2X1 _13153_ (
    .A(_05948_),
    .B(_05977_),
    .Y(_05978_)
  );
  AOI21X1 _13154_ (
    .A(_05961_),
    .B(_05975_),
    .C(_05978_),
    .Y(_05979_)
  );
  INVX1 _13155_ (
    .A(_05979_),
    .Y(_05980_)
  );
  NOR2X1 _13156_ (
    .A(_00127_),
    .B(_00128_),
    .Y(_05981_)
  );
  NOR2X1 _13157_ (
    .A(_00106_),
    .B(_00105_),
    .Y(_05982_)
  );
  NAND3X1 _13158_ (
    .A(_05926_),
    .B(_00107_),
    .C(_05982_),
    .Y(_05983_)
  );
  NOR2X1 _13159_ (
    .A(_00102_),
    .B(_00101_),
    .Y(_05984_)
  );
  NOR2X1 _13160_ (
    .A(_00103_),
    .B(_05924_),
    .Y(_05985_)
  );
  NAND2X1 _13161_ (
    .A(_05984_),
    .B(_05985_),
    .Y(_05986_)
  );
  NOR2X1 _13162_ (
    .A(_05983_),
    .B(_05986_),
    .Y(_05987_)
  );
  NAND3X1 _13163_ (
    .A(_05927_),
    .B(_00126_),
    .C(_05928_),
    .Y(_05988_)
  );
  NOR2X1 _13164_ (
    .A(_00098_),
    .B(_00109_),
    .Y(_05989_)
  );
  NOR2X1 _13165_ (
    .A(_00100_),
    .B(_00099_),
    .Y(_05990_)
  );
  NAND2X1 _13166_ (
    .A(_05989_),
    .B(_05990_),
    .Y(_05991_)
  );
  NOR2X1 _13167_ (
    .A(_05988_),
    .B(_05991_),
    .Y(_05992_)
  );
  NOR2X1 _13168_ (
    .A(_00105_),
    .B(_00108_),
    .Y(_05993_)
  );
  NOR2X1 _13169_ (
    .A(_00102_),
    .B(_05924_),
    .Y(_05994_)
  );
  OR2X1 _13170_ (
    .A(_00109_),
    .B(_00100_),
    .Y(_05995_)
  );
  NOR2X1 _13171_ (
    .A(1'h0),
    .B(_05995_),
    .Y(_05996_)
  );
  NAND3X1 _13172_ (
    .A(_05993_),
    .B(_05994_),
    .C(_05996_),
    .Y(_05997_)
  );
  NOR2X1 _13173_ (
    .A(_00101_),
    .B(_00103_),
    .Y(_05998_)
  );
  NAND3X1 _13174_ (
    .A(_05925_),
    .B(_00107_),
    .C(_05998_),
    .Y(_05999_)
  );
  NOR2X1 _13175_ (
    .A(_00098_),
    .B(_00099_),
    .Y(_06000_)
  );
  NAND3X1 _13176_ (
    .A(_00126_),
    .B(_05928_),
    .C(_06000_),
    .Y(_06001_)
  );
  OR2X1 _13177_ (
    .A(_05999_),
    .B(_06001_),
    .Y(_06002_)
  );
  NOR2X1 _13178_ (
    .A(_05997_),
    .B(_06002_),
    .Y(_06003_)
  );
  OAI21X1 _13179_ (
    .A(_00127_),
    .B(_00128_),
    .C(_06003_),
    .Y(_06004_)
  );
  NOR2X1 _13180_ (
    .A(_00114_),
    .B(_00116_),
    .Y(_06005_)
  );
  NAND2X1 _13181_ (
    .A(_00125_),
    .B(_00112_),
    .Y(_06006_)
  );
  NOR2X1 _13182_ (
    .A(_00124_),
    .B(_00111_),
    .Y(_06007_)
  );
  NAND3X1 _13183_ (
    .A(_00113_),
    .B(_00115_),
    .C(_06007_),
    .Y(_06008_)
  );
  NOR2X1 _13184_ (
    .A(_06006_),
    .B(_06008_),
    .Y(_06009_)
  );
  AOI21X1 _13185_ (
    .A(_06005_),
    .B(_06009_),
    .C(_06004_),
    .Y(_06010_)
  );
  INVX1 _13186_ (
    .A(_06010_),
    .Y(_06011_)
  );
  AOI21X1 _13187_ (
    .A(_05971_),
    .B(_05980_),
    .C(_06010_),
    .Y(_06012_)
  );
  OAI21X1 _13188_ (
    .A(_05970_),
    .B(_05979_),
    .C(_06011_),
    .Y(_06013_)
  );
  NOR2X1 _13189_ (
    .A(_05935_),
    .B(_06004_),
    .Y(_06014_)
  );
  NAND2X1 _13190_ (
    .A(watchdog_0.wdtcnt_0_ ),
    .B(_05975_),
    .Y(_06015_)
  );
  XNOR2X1 _13191_ (
    .A(watchdog_0.wdtcnt_0_ ),
    .B(_05975_),
    .Y(_06016_)
  );
  NOR3X1 _13192_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06016_),
    .Y(_05896_)
  );
  NOR2X1 _13193_ (
    .A(_05930_),
    .B(_06015_),
    .Y(_06017_)
  );
  XNOR2X1 _13194_ (
    .A(_05930_),
    .B(_06015_),
    .Y(_06018_)
  );
  NOR3X1 _13195_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06018_),
    .Y(_05903_)
  );
  AND2X1 _13196_ (
    .A(watchdog_0.wdtcnt_2_ ),
    .B(_06017_),
    .Y(_06019_)
  );
  XNOR2X1 _13197_ (
    .A(watchdog_0.wdtcnt_2_ ),
    .B(_06017_),
    .Y(_06020_)
  );
  NOR3X1 _13198_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06020_),
    .Y(_05904_)
  );
  AND2X1 _13199_ (
    .A(_05940_),
    .B(_06017_),
    .Y(_06021_)
  );
  XNOR2X1 _13200_ (
    .A(watchdog_0.wdtcnt_3_ ),
    .B(_06019_),
    .Y(_06022_)
  );
  NOR3X1 _13201_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06022_),
    .Y(_05905_)
  );
  NAND2X1 _13202_ (
    .A(watchdog_0.wdtcnt_4_ ),
    .B(_06021_),
    .Y(_06023_)
  );
  XNOR2X1 _13203_ (
    .A(watchdog_0.wdtcnt_4_ ),
    .B(_06021_),
    .Y(_06024_)
  );
  NOR3X1 _13204_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06024_),
    .Y(_05906_)
  );
  XOR2X1 _13205_ (
    .A(watchdog_0.wdtcnt_5_ ),
    .B(_06023_),
    .Y(_06025_)
  );
  NOR3X1 _13206_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06025_),
    .Y(_05907_)
  );
  AOI21X1 _13207_ (
    .A(watchdog_0.wdtcnt_6_ ),
    .B(_05976_),
    .C(_05978_),
    .Y(_06026_)
  );
  NOR3X1 _13208_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06026_),
    .Y(_05908_)
  );
  NAND2X1 _13209_ (
    .A(_05948_),
    .B(_05975_),
    .Y(_06027_)
  );
  XOR2X1 _13210_ (
    .A(watchdog_0.wdtcnt_7_ ),
    .B(_06027_),
    .Y(_06028_)
  );
  NAND3X1 _13211_ (
    .A(watchdog_0.wdtcnt_7_ ),
    .B(_05948_),
    .C(_05975_),
    .Y(_06029_)
  );
  NOR3X1 _13212_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06028_),
    .Y(_05909_)
  );
  XOR2X1 _13213_ (
    .A(watchdog_0.wdtcnt_8_ ),
    .B(_06029_),
    .Y(_06030_)
  );
  NOR3X1 _13214_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06030_),
    .Y(_05910_)
  );
  NAND3X1 _13215_ (
    .A(watchdog_0.wdtcnt_9_ ),
    .B(_05951_),
    .C(_05975_),
    .Y(_06031_)
  );
  OAI21X1 _13216_ (
    .A(_05952_),
    .B(_05976_),
    .C(_05933_),
    .Y(_06032_)
  );
  NAND2X1 _13217_ (
    .A(_06031_),
    .B(_06032_),
    .Y(_06033_)
  );
  NOR3X1 _13218_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06033_),
    .Y(_05911_)
  );
  NOR2X1 _13219_ (
    .A(_05934_),
    .B(_06031_),
    .Y(_06034_)
  );
  XNOR2X1 _13220_ (
    .A(_05934_),
    .B(_06031_),
    .Y(_06035_)
  );
  NOR3X1 _13221_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06035_),
    .Y(_05897_)
  );
  NOR2X1 _13222_ (
    .A(_05938_),
    .B(_06031_),
    .Y(_06036_)
  );
  OAI22X1 _13223_ (
    .A(_05938_),
    .B(_06031_),
    .C(_06034_),
    .D(watchdog_0.wdtcnt_11_ ),
    .Y(_06037_)
  );
  NOR3X1 _13224_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06037_),
    .Y(_05898_)
  );
  XNOR2X1 _13225_ (
    .A(watchdog_0.wdtcnt_12_ ),
    .B(_06036_),
    .Y(_06038_)
  );
  NOR3X1 _13226_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06038_),
    .Y(_05899_)
  );
  NAND2X1 _13227_ (
    .A(_05960_),
    .B(_05975_),
    .Y(_06039_)
  );
  OAI21X1 _13228_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(_05975_),
    .C(_06039_),
    .Y(_06040_)
  );
  NOR3X1 _13229_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06040_),
    .Y(_05900_)
  );
  NAND3X1 _13230_ (
    .A(watchdog_0.wdtcnt_13_ ),
    .B(_05953_),
    .C(_05975_),
    .Y(_06041_)
  );
  XOR2X1 _13231_ (
    .A(watchdog_0.wdtcnt_14_ ),
    .B(_06041_),
    .Y(_06042_)
  );
  NOR3X1 _13232_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06042_),
    .Y(_05901_)
  );
  NAND2X1 _13233_ (
    .A(_05955_),
    .B(_05975_),
    .Y(_06043_)
  );
  OAI21X1 _13234_ (
    .A(watchdog_0.wdtcnt_15_ ),
    .B(_05975_),
    .C(_06043_),
    .Y(_06044_)
  );
  NOR3X1 _13235_ (
    .A(_06013_),
    .B(_06014_),
    .C(_06044_),
    .Y(_05902_)
  );
  MUX2X1 _13236_ (
    .A(watchdog_0.wdtctl_0_ ),
    .B(_00110_),
    .S(_06004_),
    .Y(_06045_)
  );
  INVX1 _13237_ (
    .A(_06045_),
    .Y(_05912_)
  );
  MUX2X1 _13238_ (
    .A(watchdog_0.wdtctl_1_ ),
    .B(_00117_),
    .S(_06004_),
    .Y(_06046_)
  );
  INVX1 _13239_ (
    .A(_06046_),
    .Y(_05913_)
  );
  MUX2X1 _13240_ (
    .A(watchdog_0.wdtctl_2_ ),
    .B(_00118_),
    .S(_06004_),
    .Y(_06047_)
  );
  INVX1 _13241_ (
    .A(_06047_),
    .Y(_05914_)
  );
  AND2X1 _13242_ (
    .A(watchdog_0.wdtctl_3_ ),
    .B(_06004_),
    .Y(_05915_)
  );
  MUX2X1 _13243_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(_00120_),
    .S(_06004_),
    .Y(_06048_)
  );
  INVX1 _13244_ (
    .A(_06048_),
    .Y(_05916_)
  );
  AND2X1 _13245_ (
    .A(watchdog_0.wdtctl_5_ ),
    .B(_06004_),
    .Y(_05917_)
  );
  AND2X1 _13246_ (
    .A(sfr_0.UNUSED_wdtnmies ),
    .B(_06004_),
    .Y(_05918_)
  );
  MUX2X1 _13247_ (
    .A(watchdog_0.wdtctl_7_ ),
    .B(_00123_),
    .S(_06004_),
    .Y(_06049_)
  );
  INVX1 _13248_ (
    .A(_06049_),
    .Y(_05919_)
  );
  NAND2X1 _13249_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(_00084_),
    .Y(_06050_)
  );
  NAND3X1 _13250_ (
    .A(_05936_),
    .B(sfr_0.ifg1_0_ ),
    .C(_06050_),
    .Y(_06051_)
  );
  NAND3X1 _13251_ (
    .A(_05937_),
    .B(_06012_),
    .C(_06051_),
    .Y(_05920_)
  );
  NAND3X1 _13252_ (
    .A(_05981_),
    .B(_05987_),
    .C(_05992_),
    .Y(_06052_)
  );
  INVX1 _13253_ (
    .A(_06052_),
    .Y(per_dout_wdog_11_)
  );
  NAND3X1 _13254_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(sfr_0.ifg1_0_ ),
    .C(sfr_0.ie1_0_ ),
    .Y(_06053_)
  );
  INVX1 _13255_ (
    .A(_06053_),
    .Y(frontend_0.wdt_irq )
  );
  AOI22X1 _13256_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(_06011_),
    .C(_06012_),
    .D(_05937_),
    .Y(_05895_)
  );
  NOR2X1 _13257_ (
    .A(_05931_),
    .B(_06052_),
    .Y(per_dout_wdog_0_)
  );
  NOR2X1 _13258_ (
    .A(_05932_),
    .B(_06052_),
    .Y(per_dout_wdog_1_)
  );
  AND2X1 _13259_ (
    .A(watchdog_0.wdtctl_2_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_2_)
  );
  AND2X1 _13260_ (
    .A(watchdog_0.wdtctl_3_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_3_)
  );
  AND2X1 _13261_ (
    .A(watchdog_0.wdtctl_4_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_4_)
  );
  AND2X1 _13262_ (
    .A(watchdog_0.wdtctl_5_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_5_)
  );
  AND2X1 _13263_ (
    .A(sfr_0.UNUSED_wdtnmies ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_6_)
  );
  AND2X1 _13264_ (
    .A(watchdog_0.wdtctl_7_ ),
    .B(per_dout_wdog_11_),
    .Y(per_dout_wdog_7_)
  );
  DFFSR _13265_ (
    .CLK(dco_clk),
    .D(_05895_),
    .Q(clock_module_0.wdt_reset ),
    .R(_05921_),
    .S(1'h1)
  );
  DFFSR _13266_ (
    .CLK(dco_clk),
    .D(_05920_),
    .Q(sfr_0.ifg1_0_ ),
    .R(_05921_),
    .S(1'h1)
  );
  DFFSR _13267_ (
    .CLK(dco_clk),
    .D(_05896_),
    .Q(watchdog_0.wdtcnt_0_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13268_ (
    .CLK(dco_clk),
    .D(_05903_),
    .Q(watchdog_0.wdtcnt_1_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13269_ (
    .CLK(dco_clk),
    .D(_05904_),
    .Q(watchdog_0.wdtcnt_2_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13270_ (
    .CLK(dco_clk),
    .D(_05905_),
    .Q(watchdog_0.wdtcnt_3_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13271_ (
    .CLK(dco_clk),
    .D(_05906_),
    .Q(watchdog_0.wdtcnt_4_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13272_ (
    .CLK(dco_clk),
    .D(_05907_),
    .Q(watchdog_0.wdtcnt_5_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13273_ (
    .CLK(dco_clk),
    .D(_05908_),
    .Q(watchdog_0.wdtcnt_6_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13274_ (
    .CLK(dco_clk),
    .D(_05909_),
    .Q(watchdog_0.wdtcnt_7_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13275_ (
    .CLK(dco_clk),
    .D(_05910_),
    .Q(watchdog_0.wdtcnt_8_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13276_ (
    .CLK(dco_clk),
    .D(_05911_),
    .Q(watchdog_0.wdtcnt_9_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13277_ (
    .CLK(dco_clk),
    .D(_05897_),
    .Q(watchdog_0.wdtcnt_10_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13278_ (
    .CLK(dco_clk),
    .D(_05898_),
    .Q(watchdog_0.wdtcnt_11_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13279_ (
    .CLK(dco_clk),
    .D(_05899_),
    .Q(watchdog_0.wdtcnt_12_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13280_ (
    .CLK(dco_clk),
    .D(_05900_),
    .Q(watchdog_0.wdtcnt_13_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13281_ (
    .CLK(dco_clk),
    .D(_05901_),
    .Q(watchdog_0.wdtcnt_14_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13282_ (
    .CLK(dco_clk),
    .D(_05902_),
    .Q(watchdog_0.wdtcnt_15_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13283_ (
    .CLK(dco_clk),
    .D(_05912_),
    .Q(watchdog_0.wdtctl_0_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13284_ (
    .CLK(dco_clk),
    .D(_05913_),
    .Q(watchdog_0.wdtctl_1_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13285_ (
    .CLK(dco_clk),
    .D(_05914_),
    .Q(watchdog_0.wdtctl_2_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13286_ (
    .CLK(dco_clk),
    .D(_05915_),
    .Q(watchdog_0.wdtctl_3_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13287_ (
    .CLK(dco_clk),
    .D(_05916_),
    .Q(watchdog_0.wdtctl_4_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13288_ (
    .CLK(dco_clk),
    .D(_05917_),
    .Q(watchdog_0.wdtctl_5_ ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13289_ (
    .CLK(dco_clk),
    .D(_05918_),
    .Q(sfr_0.UNUSED_wdtnmies ),
    .R(_05922_),
    .S(1'h1)
  );
  DFFSR _13290_ (
    .CLK(dco_clk),
    .D(_05919_),
    .Q(watchdog_0.wdtctl_7_ ),
    .R(_05922_),
    .S(1'h1)
  );
endmodule
